* NGSPICE file created from alu.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd1_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd1_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_4 abstract view
.subckt sky130_fd_sc_hd__a2111oi_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

.subckt alu A[0] A[1] A[2] A[3] A[4] A[5] A[6] A[7] B[0] B[1] B[2] B[3] B[4] B[5]
+ B[6] B[7] VGND VPWR opcode[0] opcode[1] opcode[2] out[0] out[1] out[2] out[3] out[4]
+ out[5] out[6] out[7]
XFILLER_0_4_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_432_ _106_ net39 _108_ VGND VGND VPWR VPWR _109_ sky130_fd_sc_hd__nand3_2
X_501_ _175_ _177_ VGND VGND VPWR VPWR _178_ sky130_fd_sc_hd__nand2_1
X_294_ _219_ _222_ VGND VGND VPWR VPWR _223_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_15_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_363_ _019_ _041_ VGND VGND VPWR VPWR _042_ sky130_fd_sc_hd__and2_1
XFILLER_0_13_73 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_346_ _022_ _024_ VGND VGND VPWR VPWR _025_ sky130_fd_sc_hd__and2_2
X_415_ _090_ _091_ VGND VGND VPWR VPWR _092_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_20_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_277_ _182_ _197_ _205_ VGND VGND VPWR VPWR _207_ sky130_fd_sc_hd__and3_4
XFILLER_0_4_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_329_ _005_ _006_ _008_ VGND VGND VPWR VPWR _009_ sky130_fd_sc_hd__and3_1
XFILLER_0_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_8_Left_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_5 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_142 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput20 net20 VGND VGND VPWR VPWR out[0] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_18_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_21_Left_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_431_ _072_ _067_ _066_ VGND VGND VPWR VPWR _108_ sky130_fd_sc_hd__a21bo_1
X_362_ _021_ _040_ VGND VGND VPWR VPWR _041_ sky130_fd_sc_hd__xnor2_1
X_293_ _183_ _220_ _221_ VGND VGND VPWR VPWR _222_ sky130_fd_sc_hd__a21bo_1
X_500_ _187_ _133_ _135_ _200_ _181_ VGND VGND VPWR VPWR _177_ sky130_fd_sc_hd__o221a_1
Xrebuffer8 _075_ VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__buf_6
XFILLER_0_13_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_276_ _183_ net40 _197_ VGND VGND VPWR VPWR _206_ sky130_fd_sc_hd__a21oi_2
X_414_ _176_ net15 _089_ VGND VGND VPWR VPWR _091_ sky130_fd_sc_hd__a21oi_2
X_345_ _023_ VGND VGND VPWR VPWR _024_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_328_ net1 _218_ _221_ _007_ VGND VGND VPWR VPWR _008_ sky130_fd_sc_hd__a31o_1
XFILLER_0_10_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_259_ net19 _185_ VGND VGND VPWR VPWR _190_ sky130_fd_sc_hd__nor2_4
XPHY_EDGE_ROW_24_Left_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_73 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_95 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_6 net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_110 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput21 net21 VGND VGND VPWR VPWR out[1] sky130_fd_sc_hd__buf_2
XFILLER_0_7_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_95 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_361_ _218_ _241_ _227_ _205_ VGND VGND VPWR VPWR _040_ sky130_fd_sc_hd__o31a_1
Xrebuffer9 _075_ VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_2_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_430_ _105_ _099_ _100_ VGND VGND VPWR VPWR _107_ sky130_fd_sc_hd__nand3_2
X_292_ net2 net35 _217_ _182_ VGND VGND VPWR VPWR _221_ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_275_ net17 net18 net19 VGND VGND VPWR VPWR _205_ sky130_fd_sc_hd__nand3b_4
X_344_ net1 net2 net12 net13 VGND VGND VPWR VPWR _023_ sky130_fd_sc_hd__and4_1
X_413_ net1 net15 _089_ VGND VGND VPWR VPWR _090_ sky130_fd_sc_hd__and3_2
XFILLER_0_19_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_327_ _182_ net2 net35 _217_ VGND VGND VPWR VPWR _007_ sky130_fd_sc_hd__and4_1
X_258_ _186_ _180_ VGND VGND VPWR VPWR _189_ sky130_fd_sc_hd__nor2_4
XFILLER_0_10_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput22 net22 VGND VGND VPWR VPWR out[2] sky130_fd_sc_hd__buf_2
XFILLER_0_9_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_63 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_360_ _189_ _037_ _038_ VGND VGND VPWR VPWR _039_ sky130_fd_sc_hd__and3_1
X_291_ _193_ _197_ _217_ VGND VGND VPWR VPWR _220_ sky130_fd_sc_hd__and3_1
XFILLER_0_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_489_ _163_ _162_ _164_ VGND VGND VPWR VPWR _165_ sky130_fd_sc_hd__a21o_1
XFILLER_0_1_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_274_ net1 _183_ VGND VGND VPWR VPWR _204_ sky130_fd_sc_hd__or2b_2
X_343_ net2 net12 _021_ net1 VGND VGND VPWR VPWR _022_ sky130_fd_sc_hd__a22o_1
X_412_ net1 net14 _070_ _069_ VGND VGND VPWR VPWR _089_ sky130_fd_sc_hd__a31o_1
XFILLER_0_4_52 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_326_ _003_ _004_ _002_ VGND VGND VPWR VPWR _006_ sky130_fd_sc_hd__o21ai_2
X_257_ _176_ _183_ _187_ VGND VGND VPWR VPWR _188_ sky130_fd_sc_hd__nand3_1
XFILLER_0_10_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_309_ _217_ _195_ _226_ _237_ VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_21_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput23 net23 VGND VGND VPWR VPWR out[3] sky130_fd_sc_hd__buf_2
XFILLER_0_27_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_290_ _176_ _218_ VGND VGND VPWR VPWR _219_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_488_ _099_ _107_ VGND VGND VPWR VPWR _164_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_273_ net19 _180_ _185_ VGND VGND VPWR VPWR _203_ sky130_fd_sc_hd__and3_2
X_342_ net13 VGND VGND VPWR VPWR _021_ sky130_fd_sc_hd__buf_6
X_411_ net30 _074_ net37 VGND VGND VPWR VPWR _088_ sky130_fd_sc_hd__nand3_2
XFILLER_0_24_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_256_ net17 _186_ VGND VGND VPWR VPWR _187_ sky130_fd_sc_hd__nand2_2
XFILLER_0_19_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_325_ _002_ _003_ _004_ VGND VGND VPWR VPWR _005_ sky130_fd_sc_hd__or3_4
XFILLER_0_10_67 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_308_ _231_ _232_ _236_ _195_ VGND VGND VPWR VPWR _237_ sky130_fd_sc_hd__a211o_1
XFILLER_0_1_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput24 net24 VGND VGND VPWR VPWR out[4] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_15_Left_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_487_ _153_ _154_ _161_ VGND VGND VPWR VPWR _163_ sky130_fd_sc_hd__nand3_2
XFILLER_0_1_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_341_ _176_ _241_ _010_ _009_ VGND VGND VPWR VPWR _020_ sky130_fd_sc_hd__a31o_1
X_410_ _052_ _195_ _087_ VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__a21oi_1
X_272_ _193_ _197_ _198_ _201_ VGND VGND VPWR VPWR _202_ sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_0_Left_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_255_ net19 VGND VGND VPWR VPWR _186_ sky130_fd_sc_hd__inv_2
X_324_ _196_ net3 _238_ _182_ VGND VGND VPWR VPWR _004_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_10_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_3_Left_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_89 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_307_ _217_ _218_ _190_ _235_ VGND VGND VPWR VPWR _236_ sky130_fd_sc_hd__a31o_1
XFILLER_0_15_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput25 net25 VGND VGND VPWR VPWR out[5] sky130_fd_sc_hd__buf_2
XFILLER_0_7_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_486_ _154_ _153_ _161_ VGND VGND VPWR VPWR _162_ sky130_fd_sc_hd__a21o_1
X_271_ _193_ _197_ _200_ VGND VGND VPWR VPWR _201_ sky130_fd_sc_hd__a21oi_1
X_340_ net5 VGND VGND VPWR VPWR _019_ sky130_fd_sc_hd__buf_8
X_469_ _182_ net35 net7 net8 VGND VGND VPWR VPWR _145_ sky130_fd_sc_hd__and4_1
X_254_ net17 net18 VGND VGND VPWR VPWR _185_ sky130_fd_sc_hd__nand2_2
X_323_ net9 net10 net3 net4 VGND VGND VPWR VPWR _003_ sky130_fd_sc_hd__and4_4
XFILLER_0_27_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_167 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_24 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_306_ _217_ _218_ _198_ _234_ VGND VGND VPWR VPWR _235_ sky130_fd_sc_hd__o22a_1
XFILLER_0_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput26 net26 VGND VGND VPWR VPWR out[6] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_17_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_485_ _090_ _160_ VGND VGND VPWR VPWR _161_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_14_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_270_ _199_ VGND VGND VPWR VPWR _200_ sky130_fd_sc_hd__buf_2
XFILLER_0_24_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_468_ net35 net7 net8 _182_ VGND VGND VPWR VPWR _144_ sky130_fd_sc_hd__a22oi_2
X_399_ net29 _074_ net36 VGND VGND VPWR VPWR _077_ sky130_fd_sc_hd__a21oi_2
X_322_ net2 _218_ VGND VGND VPWR VPWR _002_ sky130_fd_sc_hd__nand2_2
XFILLER_0_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_253_ _176_ _183_ VGND VGND VPWR VPWR _184_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_305_ _200_ _233_ VGND VGND VPWR VPWR _234_ sky130_fd_sc_hd__and2b_1
Xoutput27 net27 VGND VGND VPWR VPWR out[7] sky130_fd_sc_hd__buf_8
XFILLER_0_27_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_484_ _156_ _159_ VGND VGND VPWR VPWR _160_ sky130_fd_sc_hd__xnor2_2
XPHY_EDGE_ROW_19_Left_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_467_ _218_ _238_ _021_ _052_ VGND VGND VPWR VPWR _143_ sky130_fd_sc_hd__nand4_4
X_398_ _075_ _074_ _073_ VGND VGND VPWR VPWR _076_ sky130_fd_sc_hd__and3_4
X_252_ _182_ VGND VGND VPWR VPWR _183_ sky130_fd_sc_hd__clkbuf_4
X_321_ _176_ _241_ VGND VGND VPWR VPWR _001_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_38 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_304_ net3 net11 VGND VGND VPWR VPWR _233_ sky130_fd_sc_hd__nand2_4
XFILLER_0_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_7_Left_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_158 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_483_ _157_ _158_ VGND VGND VPWR VPWR _159_ sky130_fd_sc_hd__xor2_2
XFILLER_0_24_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Left_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_466_ _238_ _021_ _052_ net11 VGND VGND VPWR VPWR _142_ sky130_fd_sc_hd__a22o_4
X_397_ _025_ _032_ _031_ VGND VGND VPWR VPWR _075_ sky130_fd_sc_hd__a21o_1
XFILLER_0_5_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_251_ net9 VGND VGND VPWR VPWR _182_ sky130_fd_sc_hd__buf_6
X_320_ _246_ _247_ _203_ VGND VGND VPWR VPWR _000_ sky130_fd_sc_hd__and3b_1
XFILLER_0_19_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_449_ net7 net15 _200_ VGND VGND VPWR VPWR _126_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_23_Left_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_303_ _229_ _230_ _203_ VGND VGND VPWR VPWR _232_ sky130_fd_sc_hd__o21a_1
XFILLER_0_1_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_482_ net2 net15 VGND VGND VPWR VPWR _158_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_20_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_396_ _072_ _066_ _067_ VGND VGND VPWR VPWR _074_ sky130_fd_sc_hd__nand3_4
X_465_ _079_ _088_ _111_ _112_ VGND VGND VPWR VPWR _141_ sky130_fd_sc_hd__a211o_4
XFILLER_0_14_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_250_ net19 _180_ VGND VGND VPWR VPWR _181_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_448_ _119_ _123_ _203_ VGND VGND VPWR VPWR _125_ sky130_fd_sc_hd__o21a_1
X_379_ _052_ _055_ VGND VGND VPWR VPWR _057_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_9_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_302_ _229_ _230_ VGND VGND VPWR VPWR _231_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_135 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_481_ net1 net16 VGND VGND VPWR VPWR _157_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_464_ _131_ _136_ _137_ _139_ _203_ VGND VGND VPWR VPWR _140_ sky130_fd_sc_hd__o311a_1
XFILLER_0_8_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_395_ _067_ _066_ _072_ VGND VGND VPWR VPWR _073_ sky130_fd_sc_hd__a21o_1
XFILLER_0_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_378_ _052_ _055_ VGND VGND VPWR VPWR _056_ sky130_fd_sc_hd__and2_1
X_447_ _119_ _123_ VGND VGND VPWR VPWR _124_ sky130_fd_sc_hd__nand2_1
X_301_ _204_ _209_ _208_ VGND VGND VPWR VPWR _230_ sky130_fd_sc_hd__a21o_1
XFILLER_0_23_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_480_ net2 net14 _103_ _155_ VGND VGND VPWR VPWR _156_ sky130_fd_sc_hd__a31o_1
XFILLER_0_0_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_463_ _119_ _123_ _138_ _130_ VGND VGND VPWR VPWR _139_ sky130_fd_sc_hd__a211o_1
X_394_ _068_ _071_ VGND VGND VPWR VPWR _072_ sky130_fd_sc_hd__xnor2_4
XTAP_TAPCELL_ROW_13_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_377_ net14 _054_ VGND VGND VPWR VPWR _055_ sky130_fd_sc_hd__xnor2_1
X_446_ _122_ net7 VGND VGND VPWR VPWR _123_ sky130_fd_sc_hd__xor2_2
XTAP_TAPCELL_ROW_0_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_9_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_300_ _217_ _228_ VGND VGND VPWR VPWR _229_ sky130_fd_sc_hd__xor2_2
XFILLER_0_15_118 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_429_ _099_ _100_ _105_ VGND VGND VPWR VPWR _106_ sky130_fd_sc_hd__a21o_1
Xinput1 A[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_27_Left_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_11_Left_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_95 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_176 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_95 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_14_Left_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_393_ _069_ _070_ VGND VGND VPWR VPWR _071_ sky130_fd_sc_hd__and2b_1
X_462_ _136_ _137_ VGND VGND VPWR VPWR _138_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_13_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_376_ _021_ _205_ _040_ VGND VGND VPWR VPWR _054_ sky130_fd_sc_hd__a21o_1
X_445_ _121_ net15 VGND VGND VPWR VPWR _122_ sky130_fd_sc_hd__xor2_2
XFILLER_0_24_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_359_ _013_ _035_ _036_ VGND VGND VPWR VPWR _038_ sky130_fd_sc_hd__nand3b_4
X_428_ _101_ _104_ VGND VGND VPWR VPWR _105_ sky130_fd_sc_hd__xor2_1
Xinput2 A[1] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_14_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_2_Left_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_461_ _135_ _132_ VGND VGND VPWR VPWR _137_ sky130_fd_sc_hd__and2b_1
X_392_ net3 net12 net13 net2 VGND VGND VPWR VPWR _070_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_444_ net41 _120_ VGND VGND VPWR VPWR _121_ sky130_fd_sc_hd__nand2_2
X_375_ _044_ _045_ _042_ VGND VGND VPWR VPWR _053_ sky130_fd_sc_hd__a21o_1
XFILLER_0_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_106 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_427_ _217_ _102_ _103_ VGND VGND VPWR VPWR _104_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_358_ _035_ _036_ _013_ VGND VGND VPWR VPWR _037_ sky130_fd_sc_hd__a21bo_1
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput3 A[2] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_289_ net11 VGND VGND VPWR VPWR _218_ sky130_fd_sc_hd__buf_8
XFILLER_0_11_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_391_ net2 net3 net12 net13 VGND VGND VPWR VPWR _069_ sky130_fd_sc_hd__and4_1
X_460_ _132_ _135_ VGND VGND VPWR VPWR _136_ sky130_fd_sc_hd__and2b_1
XFILLER_0_27_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_374_ net6 VGND VGND VPWR VPWR _052_ sky130_fd_sc_hd__buf_6
X_443_ net14 _054_ VGND VGND VPWR VPWR _120_ sky130_fd_sc_hd__or2_4
XFILLER_0_26_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput4 A[3] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__buf_4
X_288_ net3 VGND VGND VPWR VPWR _217_ sky130_fd_sc_hd__clkbuf_4
X_426_ net4 net12 _021_ net3 VGND VGND VPWR VPWR _103_ sky130_fd_sc_hd__a22o_2
X_357_ _020_ _034_ VGND VGND VPWR VPWR _036_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_409_ _203_ _059_ _086_ VGND VGND VPWR VPWR _087_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_7_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_390_ net1 net14 VGND VGND VPWR VPWR _068_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_18_Left_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_373_ _019_ _195_ _039_ _051_ VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__o2bb2a_1
X_442_ _053_ _058_ _056_ VGND VGND VPWR VPWR _119_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_287_ _193_ _195_ _202_ _216_ VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__o2bb2a_1
X_425_ _238_ net12 net13 VGND VGND VPWR VPWR _102_ sky130_fd_sc_hd__and3_1
Xinput5 A[4] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_4
X_356_ _020_ _034_ VGND VGND VPWR VPWR _035_ sky130_fd_sc_hd__nand2_2
XFILLER_0_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_408_ _189_ _081_ _082_ _085_ VGND VGND VPWR VPWR _086_ sky130_fd_sc_hd__a31o_1
XFILLER_0_7_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_55 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_339_ _238_ _195_ _000_ _018_ VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_11_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_6_Left_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_7_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_441_ _115_ _117_ VGND VGND VPWR VPWR _118_ sky130_fd_sc_hd__or2_1
X_372_ _203_ _046_ _047_ _050_ VGND VGND VPWR VPWR _051_ sky130_fd_sc_hd__a31o_1
XFILLER_0_26_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_77 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_424_ _193_ net14 VGND VGND VPWR VPWR _101_ sky130_fd_sc_hd__nand2_1
X_355_ _025_ _033_ VGND VGND VPWR VPWR _034_ sky130_fd_sc_hd__xnor2_2
X_286_ _203_ _211_ _215_ _195_ VGND VGND VPWR VPWR _216_ sky130_fd_sc_hd__a211o_1
Xinput6 A[5] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_67 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_22_Left_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_407_ _052_ net14 _190_ _194_ _084_ VGND VGND VPWR VPWR _085_ sky130_fd_sc_hd__a311o_1
X_269_ net17 net19 net18 VGND VGND VPWR VPWR _199_ sky130_fd_sc_hd__or3b_1
XFILLER_0_11_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_338_ _189_ _013_ _014_ _017_ VGND VGND VPWR VPWR _018_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_11_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_440_ _081_ _116_ _189_ VGND VGND VPWR VPWR _117_ sky130_fd_sc_hd__a21bo_1
X_371_ _019_ _021_ _190_ _194_ _049_ VGND VGND VPWR VPWR _050_ sky130_fd_sc_hd__a311o_1
XFILLER_0_25_89 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_423_ _096_ _097_ _098_ VGND VGND VPWR VPWR _100_ sky130_fd_sc_hd__a21o_1
XFILLER_0_11_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_285_ _193_ _197_ _190_ _214_ VGND VGND VPWR VPWR _215_ sky130_fd_sc_hd__a31o_1
X_354_ _031_ _032_ VGND VGND VPWR VPWR _033_ sky130_fd_sc_hd__or2b_1
Xinput7 A[6] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_1_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_268_ net18 _187_ VGND VGND VPWR VPWR _198_ sky130_fd_sc_hd__nor2_4
XFILLER_0_22_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_406_ _052_ net14 _198_ _083_ VGND VGND VPWR VPWR _084_ sky130_fd_sc_hd__o22a_1
XFILLER_0_11_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_337_ _238_ _241_ _190_ _195_ _016_ VGND VGND VPWR VPWR _017_ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_11_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput10 B[1] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_22_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_36 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_24 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_370_ _019_ _021_ _198_ _048_ VGND VGND VPWR VPWR _049_ sky130_fd_sc_hd__o22a_1
XFILLER_0_26_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_89 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_499_ net8 net16 _198_ VGND VGND VPWR VPWR _175_ sky130_fd_sc_hd__o21ai_1
X_284_ _212_ _189_ _213_ VGND VGND VPWR VPWR _214_ sky130_fd_sc_hd__and3b_1
XFILLER_0_17_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_353_ _028_ _029_ _030_ VGND VGND VPWR VPWR _032_ sky130_fd_sc_hd__a21o_1
X_422_ _096_ _097_ _098_ VGND VGND VPWR VPWR _099_ sky130_fd_sc_hd__nand3_2
XTAP_TAPCELL_ROW_1_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput8 A[7] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_2
XFILLER_0_9_130 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_14 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_267_ _196_ VGND VGND VPWR VPWR _197_ sky130_fd_sc_hd__clkbuf_4
X_336_ _238_ _241_ _198_ _015_ VGND VGND VPWR VPWR _016_ sky130_fd_sc_hd__o22a_1
X_405_ _052_ net14 _200_ VGND VGND VPWR VPWR _083_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput11 B[2] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__buf_2
X_319_ _244_ _245_ _240_ VGND VGND VPWR VPWR _247_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_22_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_48 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_112 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_36 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_498_ _172_ _173_ _189_ VGND VGND VPWR VPWR _174_ sky130_fd_sc_hd__o21a_1
XFILLER_0_5_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_421_ _062_ _061_ _060_ VGND VGND VPWR VPWR _098_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput9 B[0] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__buf_4
X_283_ _183_ _193_ _197_ _176_ VGND VGND VPWR VPWR _213_ sky130_fd_sc_hd__a22o_1
X_352_ _028_ _029_ _030_ VGND VGND VPWR VPWR _031_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_1_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_404_ _035_ _038_ _080_ VGND VGND VPWR VPWR _082_ sky130_fd_sc_hd__nand3_1
X_266_ net10 VGND VGND VPWR VPWR _196_ sky130_fd_sc_hd__buf_12
X_335_ _238_ _241_ _200_ VGND VGND VPWR VPWR _015_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput12 B[3] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_26_Left_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_249_ net17 net18 VGND VGND VPWR VPWR _180_ sky130_fd_sc_hd__or2_2
X_318_ _240_ _244_ _245_ VGND VGND VPWR VPWR _246_ sky130_fd_sc_hd__and3_1
XFILLER_0_3_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_10_Left_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Left_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_124 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_497_ _170_ _171_ net28 VGND VGND VPWR VPWR _173_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_5_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_70 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_420_ _095_ _093_ _094_ VGND VGND VPWR VPWR _097_ sky130_fd_sc_hd__nand3_2
X_351_ _002_ _004_ _003_ VGND VGND VPWR VPWR _030_ sky130_fd_sc_hd__o21bai_2
X_282_ _176_ _183_ _193_ _197_ VGND VGND VPWR VPWR _212_ sky130_fd_sc_hd__and4_1
X_403_ _035_ _038_ _080_ VGND VGND VPWR VPWR _081_ sky130_fd_sc_hd__a21o_1
X_334_ _224_ _012_ VGND VGND VPWR VPWR _014_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_176 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_265_ _194_ VGND VGND VPWR VPWR _195_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_25_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap28 _115_ VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput13 B[4] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_2
X_317_ _238_ _242_ _243_ VGND VGND VPWR VPWR _245_ sky130_fd_sc_hd__or3_2
X_248_ net1 VGND VGND VPWR VPWR _176_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_138 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_496_ _170_ net28 _171_ VGND VGND VPWR VPWR _172_ sky130_fd_sc_hd__and3_1
XFILLER_0_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_82 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_350_ _027_ net32 _233_ VGND VGND VPWR VPWR _029_ sky130_fd_sc_hd__o21ai_2
X_281_ _204_ _210_ VGND VGND VPWR VPWR _211_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_22_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_479_ net3 net4 net12 _021_ VGND VGND VPWR VPWR _155_ sky130_fd_sc_hd__and4_1
XFILLER_0_9_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_402_ _078_ net33 VGND VGND VPWR VPWR _080_ sky130_fd_sc_hd__nand2_1
X_333_ _224_ _012_ VGND VGND VPWR VPWR _013_ sky130_fd_sc_hd__nand2_2
X_264_ net19 _180_ VGND VGND VPWR VPWR _194_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput14 B[5] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_4
X_316_ _242_ _243_ _238_ VGND VGND VPWR VPWR _244_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_5_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_495_ _168_ _169_ _141_ VGND VGND VPWR VPWR _171_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_9_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_94 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_280_ _208_ _209_ VGND VGND VPWR VPWR _210_ sky130_fd_sc_hd__or2b_1
XFILLER_0_22_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_478_ _152_ _148_ _149_ VGND VGND VPWR VPWR _154_ sky130_fd_sc_hd__nand3_2
XFILLER_0_13_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_263_ net2 VGND VGND VPWR VPWR _193_ sky130_fd_sc_hd__buf_2
XFILLER_0_2_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_401_ _024_ _077_ _076_ VGND VGND VPWR VPWR _079_ sky130_fd_sc_hd__or3_4
X_332_ _001_ _011_ VGND VGND VPWR VPWR _012_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_6_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput15 B[6] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_4
X_315_ _183_ _197_ _218_ _241_ _205_ VGND VGND VPWR VPWR _243_ sky130_fd_sc_hd__o311a_1
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_494_ _169_ _168_ _141_ VGND VGND VPWR VPWR _170_ sky130_fd_sc_hd__or3_4
XFILLER_0_10_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_17_Left_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_477_ _149_ _148_ _152_ VGND VGND VPWR VPWR _153_ sky130_fd_sc_hd__a21o_1
XFILLER_0_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_331_ _009_ _010_ VGND VGND VPWR VPWR _011_ sky130_fd_sc_hd__and2b_1
X_400_ _076_ _077_ _024_ VGND VGND VPWR VPWR _078_ sky130_fd_sc_hd__o21ai_1
X_262_ _176_ _181_ _184_ _192_ VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput16 B[7] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_2
X_314_ _218_ net40 _227_ _241_ VGND VGND VPWR VPWR _242_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_2_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Left_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_493_ _165_ _167_ _166_ VGND VGND VPWR VPWR _169_ sky130_fd_sc_hd__and3_1
X_476_ _150_ _151_ VGND VGND VPWR VPWR _152_ sky130_fd_sc_hd__xor2_2
XFILLER_0_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_330_ _005_ _006_ _008_ VGND VGND VPWR VPWR _010_ sky130_fd_sc_hd__a21o_1
X_261_ _180_ _185_ _188_ _191_ VGND VGND VPWR VPWR _192_ sky130_fd_sc_hd__a31o_1
X_459_ _133_ _134_ VGND VGND VPWR VPWR _135_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput17 opcode[0] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__buf_2
X_313_ net12 VGND VGND VPWR VPWR _241_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_492_ _165_ _166_ _167_ VGND VGND VPWR VPWR _168_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_8_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_475_ _217_ net14 VGND VGND VPWR VPWR _151_ sky130_fd_sc_hd__nand2_1
X_260_ _189_ _190_ _176_ _183_ VGND VGND VPWR VPWR _191_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_19_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_389_ _063_ _064_ _065_ VGND VGND VPWR VPWR _067_ sky130_fd_sc_hd__a21o_4
X_458_ net8 net16 VGND VGND VPWR VPWR _134_ sky130_fd_sc_hd__or2_1
X_312_ _229_ _230_ _239_ VGND VGND VPWR VPWR _240_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_16_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput18 opcode[1] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_21_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_491_ _092_ _110_ _109_ VGND VGND VPWR VPWR _167_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_19_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_474_ _095_ _094_ _093_ VGND VGND VPWR VPWR _150_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_26_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_457_ net8 net16 VGND VGND VPWR VPWR _133_ sky130_fd_sc_hd__nand2_1
X_388_ net38 _064_ _065_ VGND VGND VPWR VPWR _066_ sky130_fd_sc_hd__nand3_4
XTAP_TAPCELL_ROW_24_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput19 opcode[2] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__clkbuf_4
X_311_ _217_ _228_ VGND VGND VPWR VPWR _239_ sky130_fd_sc_hd__and2_1
XFILLER_0_5_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_54 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_9_Left_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_490_ _164_ _162_ _163_ VGND VGND VPWR VPWR _166_ sky130_fd_sc_hd__nand3_1
XFILLER_0_25_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_473_ _241_ _019_ _146_ _147_ VGND VGND VPWR VPWR _149_ sky130_fd_sc_hd__nand4_2
XFILLER_0_26_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_456_ net15 _120_ _205_ VGND VGND VPWR VPWR _132_ sky130_fd_sc_hd__o21ai_2
X_387_ _233_ _027_ net31 VGND VGND VPWR VPWR _065_ sky130_fd_sc_hd__o21bai_4
XFILLER_0_12_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_310_ net4 VGND VGND VPWR VPWR _238_ sky130_fd_sc_hd__buf_12
XFILLER_0_5_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_439_ net34 _114_ VGND VGND VPWR VPWR _116_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_21_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_25_Left_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_140 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_12_Left_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_472_ _241_ _019_ _146_ _147_ VGND VGND VPWR VPWR _148_ sky130_fd_sc_hd__a22o_4
XFILLER_0_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_118 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer10 _063_ VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__buf_2
XFILLER_0_6_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_455_ _119_ _123_ _130_ VGND VGND VPWR VPWR _131_ sky130_fd_sc_hd__a21oi_2
X_386_ _062_ _060_ _061_ VGND VGND VPWR VPWR _064_ sky130_fd_sc_hd__nand3_2
XFILLER_0_10_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_438_ _035_ _038_ _080_ _113_ _114_ VGND VGND VPWR VPWR _115_ sky130_fd_sc_hd__a2111oi_4
X_369_ _019_ _021_ _200_ VGND VGND VPWR VPWR _048_ sky130_fd_sc_hd__a21oi_1
Xrebuffer1 _073_ VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_471_ _144_ _145_ _142_ _143_ VGND VGND VPWR VPWR _147_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrebuffer11 _107_ VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__buf_6
XFILLER_0_13_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_454_ net7 _122_ VGND VGND VPWR VPWR _130_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_27_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_47 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_385_ _060_ _061_ _062_ VGND VGND VPWR VPWR _063_ sky130_fd_sc_hd__a21o_1
XFILLER_0_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_368_ _044_ _045_ VGND VGND VPWR VPWR _047_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_299_ _218_ _227_ VGND VGND VPWR VPWR _228_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_2_103 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer2 net29 VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__dlygate4sd1_1
X_437_ _111_ _112_ _088_ _079_ VGND VGND VPWR VPWR _114_ sky130_fd_sc_hd__o211a_1
XFILLER_0_1_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_8_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclone7 net10 VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__clkbuf_16
XFILLER_0_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_470_ _143_ _142_ _144_ _145_ VGND VGND VPWR VPWR _146_ sky130_fd_sc_hd__a211o_4
Xrebuffer12 _205_ VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__buf_2
XFILLER_0_21_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_453_ net7 _195_ _118_ _129_ VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__a22oi_2
X_384_ net11 net4 VGND VGND VPWR VPWR _062_ sky130_fd_sc_hd__and2_4
XFILLER_0_12_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_107 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_298_ _183_ _197_ _205_ VGND VGND VPWR VPWR _227_ sky130_fd_sc_hd__o21a_2
X_436_ _088_ net33 _111_ _112_ VGND VGND VPWR VPWR _113_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_2_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_367_ _044_ _045_ VGND VGND VPWR VPWR _046_ sky130_fd_sc_hd__nand2_1
Xrebuffer3 _026_ VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_419_ _093_ _094_ _095_ VGND VGND VPWR VPWR _096_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_8_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_5_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_1 _125_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_16_Left_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer13 _205_ VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__dlygate4sd1_1
X_452_ _124_ _125_ _128_ VGND VGND VPWR VPWR _129_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_27_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_383_ _196_ net5 net6 net9 VGND VGND VPWR VPWR _061_ sky130_fd_sc_hd__a22o_4
XFILLER_0_8_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_1_Left_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_366_ _240_ _245_ _244_ VGND VGND VPWR VPWR _045_ sky130_fd_sc_hd__a21bo_1
X_435_ _109_ _110_ _092_ VGND VGND VPWR VPWR _112_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_2_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_297_ _224_ _225_ VGND VGND VPWR VPWR _226_ sky130_fd_sc_hd__nor2_1
Xrebuffer4 _026_ VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_3_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_418_ net11 _019_ VGND VGND VPWR VPWR _095_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_8_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_349_ _233_ _027_ _026_ VGND VGND VPWR VPWR _028_ sky130_fd_sc_hd__or3_4
XPHY_EDGE_ROW_4_Left_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_36 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_2 _154_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_27_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_382_ _182_ _196_ _019_ net6 VGND VGND VPWR VPWR _060_ sky130_fd_sc_hd__nand4_4
X_451_ net7 net15 _190_ _195_ _127_ VGND VGND VPWR VPWR _128_ sky130_fd_sc_hd__a311o_1
X_503_ _140_ _178_ _174_ _181_ _179_ VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__o32a_4
X_296_ _212_ _223_ _189_ VGND VGND VPWR VPWR _225_ sky130_fd_sc_hd__o21ai_1
X_434_ _092_ _109_ _110_ VGND VGND VPWR VPWR _111_ sky130_fd_sc_hd__and3_4
XTAP_TAPCELL_ROW_15_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_365_ _042_ _043_ VGND VGND VPWR VPWR _044_ sky130_fd_sc_hd__nor2_1
Xrebuffer5 _079_ VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_12_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_348_ net10 net4 net5 net9 VGND VGND VPWR VPWR _027_ sky130_fd_sc_hd__a22oi_4
X_279_ _193_ _206_ _207_ VGND VGND VPWR VPWR _209_ sky130_fd_sc_hd__or3_4
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_417_ _196_ _052_ net7 _182_ VGND VGND VPWR VPWR _094_ sky130_fd_sc_hd__a22o_4
XFILLER_0_24_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_3 _246_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_381_ _053_ _058_ VGND VGND VPWR VPWR _059_ sky130_fd_sc_hd__xor2_1
X_450_ net7 net15 _198_ _126_ VGND VGND VPWR VPWR _127_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_2_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_433_ _106_ _107_ _108_ VGND VGND VPWR VPWR _110_ sky130_fd_sc_hd__a21o_2
X_502_ net8 VGND VGND VPWR VPWR _179_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_15_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_170 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrebuffer6 _113_ VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_1
X_364_ _019_ _041_ VGND VGND VPWR VPWR _043_ sky130_fd_sc_hd__nor2_1
X_295_ _212_ _223_ VGND VGND VPWR VPWR _224_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_12_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_278_ _206_ _207_ _193_ VGND VGND VPWR VPWR _208_ sky130_fd_sc_hd__o21a_1
X_416_ _182_ net35 _052_ net7 VGND VGND VPWR VPWR _093_ sky130_fd_sc_hd__nand4_4
X_347_ net4 net10 net9 net5 VGND VGND VPWR VPWR _026_ sky130_fd_sc_hd__and4_1
XFILLER_0_20_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_95 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_4 net20 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_130 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_380_ _056_ _057_ VGND VGND VPWR VPWR _058_ sky130_fd_sc_hd__nor2_2
XFILLER_0_12_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_138 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
.ends

