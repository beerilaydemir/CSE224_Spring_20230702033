VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ZeroToFiveCounter
  CLASS BLOCK ;
  FOREIGN ZeroToFiveCounter ;
  ORIGIN 0.000 0.000 ;
  SIZE 74.435 BY 85.155 ;
  PIN AN[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END AN[0]
  PIN AN[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END AN[1]
  PIN AN[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.435 64.640 74.435 65.240 ;
    END
  END AN[2]
  PIN AN[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.435 17.040 74.435 17.640 ;
    END
  END AN[3]
  PIN AN[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END AN[4]
  PIN AN[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END AN[5]
  PIN AN[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.435 68.040 74.435 68.640 ;
    END
  END AN[6]
  PIN AN[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.435 13.640 74.435 14.240 ;
    END
  END AN[7]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 15.895 10.640 17.495 73.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 31.650 10.640 33.250 73.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 47.405 10.640 49.005 73.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 63.160 10.640 64.760 73.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 21.195 68.780 22.795 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 36.830 68.780 38.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 52.465 68.780 54.065 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 68.100 68.780 69.700 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 12.595 10.640 14.195 73.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 28.350 10.640 29.950 73.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 44.105 10.640 45.705 73.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 59.860 10.640 61.460 73.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 17.895 68.780 19.495 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 33.530 68.780 35.130 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 49.165 68.780 50.765 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 64.800 68.780 66.400 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END clk
  PIN count[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END count[0]
  PIN count[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END count[1]
  PIN count[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END count[2]
  PIN count[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 70.435 20.440 74.435 21.040 ;
    END
  END count[3]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END rst
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 68.730 73.630 ;
      LAYER li1 ;
        RECT 5.520 10.795 68.540 73.525 ;
      LAYER met1 ;
        RECT 4.210 10.640 68.540 73.680 ;
      LAYER met2 ;
        RECT 4.230 4.280 67.070 73.625 ;
        RECT 4.230 4.000 35.230 4.280 ;
        RECT 36.070 4.000 44.890 4.280 ;
        RECT 45.730 4.000 48.110 4.280 ;
        RECT 48.950 4.000 51.330 4.280 ;
        RECT 52.170 4.000 67.070 4.280 ;
      LAYER met3 ;
        RECT 3.990 69.040 70.435 73.605 ;
        RECT 4.400 67.640 70.035 69.040 ;
        RECT 3.990 65.640 70.435 67.640 ;
        RECT 4.400 64.240 70.035 65.640 ;
        RECT 3.990 62.240 70.435 64.240 ;
        RECT 4.400 60.840 70.435 62.240 ;
        RECT 3.990 21.440 70.435 60.840 ;
        RECT 3.990 20.040 70.035 21.440 ;
        RECT 3.990 18.040 70.435 20.040 ;
        RECT 4.400 16.640 70.035 18.040 ;
        RECT 3.990 14.640 70.435 16.640 ;
        RECT 4.400 13.240 70.035 14.640 ;
        RECT 3.990 10.715 70.435 13.240 ;
      LAYER met4 ;
        RECT 30.655 47.775 30.985 61.705 ;
  END
END ZeroToFiveCounter
END LIBRARY

