magic
tech sky130A
magscale 1 2
timestamp 1746885429
<< checkpaint >>
rect -3932 -3932 23932 23932
<< viali >>
rect 9045 17289 9079 17323
rect 17877 17289 17911 17323
rect 2421 17221 2455 17255
rect 3893 17221 3927 17255
rect 4261 17221 4295 17255
rect 6469 17221 6503 17255
rect 9597 17221 9631 17255
rect 9781 17221 9815 17255
rect 2237 17153 2271 17187
rect 5457 17153 5491 17187
rect 9229 17153 9263 17187
rect 9413 17153 9447 17187
rect 11069 17153 11103 17187
rect 11805 17153 11839 17187
rect 14105 17153 14139 17187
rect 16405 17153 16439 17187
rect 17325 17153 17359 17187
rect 17693 17153 17727 17187
rect 18521 17153 18555 17187
rect 5365 17085 5399 17119
rect 11897 17085 11931 17119
rect 12633 17085 12667 17119
rect 16037 17085 16071 17119
rect 18245 17085 18279 17119
rect 5825 17017 5859 17051
rect 1777 16949 1811 16983
rect 2145 16949 2179 16983
rect 2513 16949 2547 16983
rect 6561 16949 6595 16983
rect 11253 16949 11287 16983
rect 14289 16949 14323 16983
rect 16589 16745 16623 16779
rect 10701 16677 10735 16711
rect 14841 16677 14875 16711
rect 16773 16677 16807 16711
rect 16865 16677 16899 16711
rect 2237 16609 2271 16643
rect 10977 16609 11011 16643
rect 11345 16609 11379 16643
rect 15209 16609 15243 16643
rect 2053 16541 2087 16575
rect 10425 16541 10459 16575
rect 11161 16541 11195 16575
rect 15117 16541 15151 16575
rect 16865 16541 16899 16575
rect 17049 16541 17083 16575
rect 17141 16541 17175 16575
rect 18245 16541 18279 16575
rect 1501 16473 1535 16507
rect 1869 16473 1903 16507
rect 10701 16473 10735 16507
rect 14565 16473 14599 16507
rect 16405 16473 16439 16507
rect 10517 16405 10551 16439
rect 16605 16405 16639 16439
rect 17877 16405 17911 16439
rect 18429 16405 18463 16439
rect 3065 16201 3099 16235
rect 16957 16201 16991 16235
rect 12725 16133 12759 16167
rect 3065 16065 3099 16099
rect 6561 16065 6595 16099
rect 6653 16065 6687 16099
rect 7021 16065 7055 16099
rect 12173 16065 12207 16099
rect 12357 16065 12391 16099
rect 12633 16065 12667 16099
rect 12909 16065 12943 16099
rect 2697 15997 2731 16031
rect 3249 15997 3283 16031
rect 6929 15861 6963 15895
rect 12265 15861 12299 15895
rect 12909 15861 12943 15895
rect 5457 15657 5491 15691
rect 8585 15657 8619 15691
rect 9505 15657 9539 15691
rect 10609 15657 10643 15691
rect 8769 15589 8803 15623
rect 14841 15589 14875 15623
rect 4721 15521 4755 15555
rect 7481 15521 7515 15555
rect 12633 15521 12667 15555
rect 3985 15453 4019 15487
rect 4169 15453 4203 15487
rect 4261 15453 4295 15487
rect 4629 15453 4663 15487
rect 5181 15453 5215 15487
rect 5273 15453 5307 15487
rect 6929 15453 6963 15487
rect 7757 15453 7791 15487
rect 8033 15453 8067 15487
rect 8309 15453 8343 15487
rect 8953 15453 8987 15487
rect 9045 15453 9079 15487
rect 9229 15453 9263 15487
rect 9321 15453 9355 15487
rect 10609 15453 10643 15487
rect 11069 15453 11103 15487
rect 11437 15453 11471 15487
rect 11713 15453 11747 15487
rect 12541 15453 12575 15487
rect 12817 15453 12851 15487
rect 13369 15453 13403 15487
rect 15025 15453 15059 15487
rect 15301 15453 15335 15487
rect 6561 15385 6595 15419
rect 7941 15385 7975 15419
rect 8401 15385 8435 15419
rect 12449 15385 12483 15419
rect 3801 15317 3835 15351
rect 4997 15317 5031 15351
rect 8601 15317 8635 15351
rect 13185 15317 13219 15351
rect 15209 15317 15243 15351
rect 1777 15113 1811 15147
rect 5273 15045 5307 15079
rect 11897 15045 11931 15079
rect 1593 14977 1627 15011
rect 1869 14977 1903 15011
rect 4537 14977 4571 15011
rect 4629 14977 4663 15011
rect 4813 14977 4847 15011
rect 9597 14977 9631 15011
rect 10149 14977 10183 15011
rect 10793 14977 10827 15011
rect 11713 14977 11747 15011
rect 12357 14977 12391 15011
rect 12541 14977 12575 15011
rect 12909 14977 12943 15011
rect 13001 14977 13035 15011
rect 13277 14977 13311 15011
rect 13369 14977 13403 15011
rect 13553 14977 13587 15011
rect 13921 14977 13955 15011
rect 14114 14977 14148 15011
rect 16681 14977 16715 15011
rect 17141 14977 17175 15011
rect 17417 14977 17451 15011
rect 18153 14977 18187 15011
rect 9689 14909 9723 14943
rect 10333 14909 10367 14943
rect 10701 14909 10735 14943
rect 14749 14909 14783 14943
rect 17601 14909 17635 14943
rect 1409 14841 1443 14875
rect 12909 14841 12943 14875
rect 10977 14773 11011 14807
rect 11529 14773 11563 14807
rect 1777 14569 1811 14603
rect 9597 14569 9631 14603
rect 16405 14569 16439 14603
rect 16957 14501 16991 14535
rect 17693 14501 17727 14535
rect 2053 14433 2087 14467
rect 2237 14433 2271 14467
rect 9229 14433 9263 14467
rect 1961 14365 1995 14399
rect 2145 14365 2179 14399
rect 4721 14365 4755 14399
rect 4997 14365 5031 14399
rect 11713 14365 11747 14399
rect 12081 14365 12115 14399
rect 13185 14365 13219 14399
rect 13369 14365 13403 14399
rect 14105 14365 14139 14399
rect 14289 14365 14323 14399
rect 14565 14365 14599 14399
rect 16129 14365 16163 14399
rect 16681 14365 16715 14399
rect 16773 14365 16807 14399
rect 9597 14297 9631 14331
rect 11897 14297 11931 14331
rect 13093 14297 13127 14331
rect 14197 14297 14231 14331
rect 16589 14297 16623 14331
rect 16957 14297 16991 14331
rect 18061 14297 18095 14331
rect 4905 14229 4939 14263
rect 9781 14229 9815 14263
rect 11345 14229 11379 14263
rect 11529 14229 11563 14263
rect 11621 14229 11655 14263
rect 13369 14229 13403 14263
rect 16405 14229 16439 14263
rect 17601 14229 17635 14263
rect 7481 14025 7515 14059
rect 8585 14025 8619 14059
rect 9229 14025 9263 14059
rect 5273 13957 5307 13991
rect 7297 13957 7331 13991
rect 7665 13957 7699 13991
rect 18429 13957 18463 13991
rect 1501 13889 1535 13923
rect 2717 13889 2751 13923
rect 2881 13889 2915 13923
rect 2973 13889 3007 13923
rect 3065 13889 3099 13923
rect 5917 13889 5951 13923
rect 6101 13889 6135 13923
rect 6377 13889 6411 13923
rect 6469 13889 6503 13923
rect 6653 13889 6687 13923
rect 6837 13889 6871 13923
rect 7849 13889 7883 13923
rect 8769 13889 8803 13923
rect 8861 13889 8895 13923
rect 8953 13889 8987 13923
rect 12173 13889 12207 13923
rect 12357 13889 12391 13923
rect 12633 13889 12667 13923
rect 13001 13889 13035 13923
rect 18061 13889 18095 13923
rect 18245 13889 18279 13923
rect 1777 13821 1811 13855
rect 5641 13821 5675 13855
rect 6193 13821 6227 13855
rect 8585 13821 8619 13855
rect 9229 13813 9263 13847
rect 3249 13685 3283 13719
rect 5089 13685 5123 13719
rect 5273 13685 5307 13719
rect 5733 13685 5767 13719
rect 7205 13685 7239 13719
rect 9045 13685 9079 13719
rect 12633 13685 12667 13719
rect 3157 13481 3191 13515
rect 5181 13481 5215 13515
rect 9505 13481 9539 13515
rect 18429 13481 18463 13515
rect 12633 13413 12667 13447
rect 5733 13345 5767 13379
rect 7113 13345 7147 13379
rect 7573 13345 7607 13379
rect 11161 13345 11195 13379
rect 2513 13277 2547 13311
rect 2605 13277 2639 13311
rect 2881 13277 2915 13311
rect 2973 13277 3007 13311
rect 3065 13277 3099 13311
rect 3249 13277 3283 13311
rect 5273 13277 5307 13311
rect 6009 13277 6043 13311
rect 6285 13277 6319 13311
rect 7021 13277 7055 13311
rect 7389 13277 7423 13311
rect 9689 13277 9723 13311
rect 9965 13277 9999 13311
rect 11253 13277 11287 13311
rect 12633 13277 12667 13311
rect 12817 13277 12851 13311
rect 12909 13277 12943 13311
rect 15117 13277 15151 13311
rect 15301 13277 15335 13311
rect 15485 13277 15519 13311
rect 18061 13277 18095 13311
rect 18245 13277 18279 13311
rect 2697 13209 2731 13243
rect 8033 13209 8067 13243
rect 9781 13209 9815 13243
rect 17049 13209 17083 13243
rect 2329 13141 2363 13175
rect 11621 13141 11655 13175
rect 6469 12937 6503 12971
rect 7573 12937 7607 12971
rect 7757 12937 7791 12971
rect 12817 12937 12851 12971
rect 3341 12869 3375 12903
rect 3433 12869 3467 12903
rect 4169 12869 4203 12903
rect 4997 12869 5031 12903
rect 9873 12869 9907 12903
rect 18429 12869 18463 12903
rect 2605 12801 2639 12835
rect 3065 12801 3099 12835
rect 3249 12801 3283 12835
rect 3709 12801 3743 12835
rect 4629 12801 4663 12835
rect 5181 12801 5215 12835
rect 5365 12801 5399 12835
rect 5457 12801 5491 12835
rect 6653 12801 6687 12835
rect 6745 12801 6779 12835
rect 7021 12801 7055 12835
rect 7576 12801 7610 12835
rect 10057 12801 10091 12835
rect 10793 12801 10827 12835
rect 10977 12801 11011 12835
rect 11069 12801 11103 12835
rect 11529 12801 11563 12835
rect 11989 12801 12023 12835
rect 12357 12801 12391 12835
rect 12633 12801 12667 12835
rect 16037 12801 16071 12835
rect 16129 12801 16163 12835
rect 16221 12801 16255 12835
rect 17325 12801 17359 12835
rect 17693 12801 17727 12835
rect 18061 12801 18095 12835
rect 2513 12733 2547 12767
rect 2973 12733 3007 12767
rect 4537 12733 4571 12767
rect 7113 12733 7147 12767
rect 10149 12733 10183 12767
rect 10517 12733 10551 12767
rect 11897 12733 11931 12767
rect 12173 12733 12207 12767
rect 16313 12733 16347 12767
rect 4813 12665 4847 12699
rect 10609 12665 10643 12699
rect 12449 12665 12483 12699
rect 12541 12665 12575 12699
rect 2329 12597 2363 12631
rect 3617 12597 3651 12631
rect 3893 12597 3927 12631
rect 6929 12597 6963 12631
rect 7205 12597 7239 12631
rect 16497 12597 16531 12631
rect 9321 12393 9355 12427
rect 10701 12393 10735 12427
rect 12725 12393 12759 12427
rect 16129 12393 16163 12427
rect 16865 12393 16899 12427
rect 17877 12393 17911 12427
rect 4353 12325 4387 12359
rect 13277 12325 13311 12359
rect 16405 12325 16439 12359
rect 3801 12257 3835 12291
rect 5917 12257 5951 12291
rect 17417 12257 17451 12291
rect 2421 12189 2455 12223
rect 3985 12189 4019 12223
rect 4261 12189 4295 12223
rect 5365 12189 5399 12223
rect 9229 12189 9263 12223
rect 10609 12189 10643 12223
rect 10793 12189 10827 12223
rect 12909 12189 12943 12223
rect 13001 12189 13035 12223
rect 13185 12189 13219 12223
rect 13461 12189 13495 12223
rect 14473 12189 14507 12223
rect 14657 12189 14691 12223
rect 16313 12189 16347 12223
rect 16497 12189 16531 12223
rect 16589 12189 16623 12223
rect 16773 12189 16807 12223
rect 17049 12189 17083 12223
rect 17141 12189 17175 12223
rect 17509 12189 17543 12223
rect 17785 12189 17819 12223
rect 18061 12189 18095 12223
rect 18153 12189 18187 12223
rect 18521 12189 18555 12223
rect 2973 12121 3007 12155
rect 4629 12121 4663 12155
rect 12357 12121 12391 12155
rect 12541 12121 12575 12155
rect 14105 12121 14139 12155
rect 14197 12121 14231 12155
rect 1961 11849 1995 11883
rect 7389 11849 7423 11883
rect 7481 11849 7515 11883
rect 1593 11781 1627 11815
rect 1809 11781 1843 11815
rect 10977 11781 11011 11815
rect 18245 11781 18279 11815
rect 3065 11713 3099 11747
rect 4905 11713 4939 11747
rect 5181 11713 5215 11747
rect 6653 11713 6687 11747
rect 6745 11713 6779 11747
rect 6837 11713 6871 11747
rect 7021 11713 7055 11747
rect 7205 11713 7239 11747
rect 7573 11713 7607 11747
rect 7757 11713 7791 11747
rect 9597 11713 9631 11747
rect 9781 11713 9815 11747
rect 11161 11713 11195 11747
rect 11253 11713 11287 11747
rect 13921 11713 13955 11747
rect 14565 11713 14599 11747
rect 17417 11713 17451 11747
rect 17601 11713 17635 11747
rect 17785 11713 17819 11747
rect 3525 11645 3559 11679
rect 5641 11645 5675 11679
rect 8033 11645 8067 11679
rect 8125 11645 8159 11679
rect 8493 11645 8527 11679
rect 13829 11645 13863 11679
rect 14381 11645 14415 11679
rect 14473 11645 14507 11679
rect 14657 11645 14691 11679
rect 4997 11577 5031 11611
rect 9689 11577 9723 11611
rect 11069 11577 11103 11611
rect 1777 11509 1811 11543
rect 6377 11509 6411 11543
rect 7849 11509 7883 11543
rect 13553 11509 13587 11543
rect 14197 11509 14231 11543
rect 4721 11305 4755 11339
rect 5549 11305 5583 11339
rect 6101 11305 6135 11339
rect 7665 11237 7699 11271
rect 15853 11237 15887 11271
rect 16405 11237 16439 11271
rect 5273 11169 5307 11203
rect 7297 11169 7331 11203
rect 7757 11169 7791 11203
rect 10149 11169 10183 11203
rect 10609 11169 10643 11203
rect 16865 11169 16899 11203
rect 1409 11101 1443 11135
rect 3985 11101 4019 11135
rect 4537 11101 4571 11135
rect 5089 11101 5123 11135
rect 5365 11101 5399 11135
rect 6009 11101 6043 11135
rect 6201 11101 6235 11135
rect 10057 11101 10091 11135
rect 10793 11101 10827 11135
rect 10977 11101 11011 11135
rect 11069 11101 11103 11135
rect 16221 11101 16255 11135
rect 16681 11101 16715 11135
rect 17049 11101 17083 11135
rect 17509 11101 17543 11135
rect 17785 11101 17819 11135
rect 18153 11101 18187 11135
rect 1685 11033 1719 11067
rect 9229 11033 9263 11067
rect 4445 10761 4479 10795
rect 13737 10761 13771 10795
rect 15301 10761 15335 10795
rect 17667 10761 17701 10795
rect 17877 10693 17911 10727
rect 17969 10693 18003 10727
rect 3065 10625 3099 10659
rect 3985 10625 4019 10659
rect 4448 10625 4482 10659
rect 5733 10625 5767 10659
rect 5825 10625 5859 10659
rect 6377 10625 6411 10659
rect 6745 10625 6779 10659
rect 6929 10625 6963 10659
rect 7205 10625 7239 10659
rect 7297 10625 7331 10659
rect 11621 10625 11655 10659
rect 11805 10625 11839 10659
rect 13277 10625 13311 10659
rect 13461 10625 13495 10659
rect 13921 10625 13955 10659
rect 14013 10625 14047 10659
rect 14105 10625 14139 10659
rect 14289 10625 14323 10659
rect 15025 10625 15059 10659
rect 15117 10625 15151 10659
rect 15399 10625 15433 10659
rect 16129 10625 16163 10659
rect 16313 10625 16347 10659
rect 16405 10625 16439 10659
rect 16773 10625 16807 10659
rect 18337 10625 18371 10659
rect 3341 10557 3375 10591
rect 5365 10557 5399 10591
rect 5457 10557 5491 10591
rect 13185 10557 13219 10591
rect 14657 10557 14691 10591
rect 15485 10557 15519 10591
rect 18153 10557 18187 10591
rect 3617 10489 3651 10523
rect 4629 10489 4663 10523
rect 6009 10489 6043 10523
rect 6653 10489 6687 10523
rect 11621 10489 11655 10523
rect 15761 10489 15795 10523
rect 17509 10489 17543 10523
rect 3433 10421 3467 10455
rect 4077 10421 4111 10455
rect 6469 10421 6503 10455
rect 15393 10421 15427 10455
rect 15945 10421 15979 10455
rect 16865 10421 16899 10455
rect 17233 10421 17267 10455
rect 17693 10421 17727 10455
rect 18061 10421 18095 10455
rect 4077 10217 4111 10251
rect 18153 10217 18187 10251
rect 7113 10149 7147 10183
rect 16037 10149 16071 10183
rect 1961 10081 1995 10115
rect 7481 10081 7515 10115
rect 17417 10081 17451 10115
rect 18317 10081 18351 10115
rect 2789 10013 2823 10047
rect 3065 10013 3099 10047
rect 3341 10013 3375 10047
rect 3525 10013 3559 10047
rect 3985 10013 4019 10047
rect 4261 10013 4295 10047
rect 7297 10013 7331 10047
rect 7573 10013 7607 10047
rect 7665 10013 7699 10047
rect 7861 10013 7895 10047
rect 16405 10013 16439 10047
rect 17049 10013 17083 10047
rect 17509 10013 17543 10047
rect 17601 10013 17635 10047
rect 17877 10013 17911 10047
rect 17969 10013 18003 10047
rect 18521 10013 18555 10047
rect 3433 9945 3467 9979
rect 17785 9945 17819 9979
rect 18245 9945 18279 9979
rect 18429 9877 18463 9911
rect 12265 9673 12299 9707
rect 2881 9605 2915 9639
rect 4813 9605 4847 9639
rect 14841 9605 14875 9639
rect 16957 9605 16991 9639
rect 1777 9537 1811 9571
rect 1869 9537 1903 9571
rect 2053 9537 2087 9571
rect 2513 9537 2547 9571
rect 3065 9537 3099 9571
rect 4629 9537 4663 9571
rect 4905 9537 4939 9571
rect 7113 9537 7147 9571
rect 7205 9537 7239 9571
rect 7757 9537 7791 9571
rect 9597 9537 9631 9571
rect 9965 9537 9999 9571
rect 10333 9537 10367 9571
rect 12173 9537 12207 9571
rect 13921 9537 13955 9571
rect 14013 9537 14047 9571
rect 14197 9537 14231 9571
rect 14657 9537 14691 9571
rect 14933 9537 14967 9571
rect 16681 9537 16715 9571
rect 16792 9537 16826 9571
rect 17233 9537 17267 9571
rect 17785 9537 17819 9571
rect 18153 9537 18187 9571
rect 3341 9469 3375 9503
rect 3801 9469 3835 9503
rect 4445 9469 4479 9503
rect 7573 9469 7607 9503
rect 8953 9469 8987 9503
rect 9689 9469 9723 9503
rect 9873 9469 9907 9503
rect 10885 9469 10919 9503
rect 17417 9469 17451 9503
rect 3249 9401 3283 9435
rect 14473 9401 14507 9435
rect 2053 9333 2087 9367
rect 2697 9333 2731 9367
rect 4261 9333 4295 9367
rect 14381 9333 14415 9367
rect 16681 9333 16715 9367
rect 1409 9129 1443 9163
rect 2697 9129 2731 9163
rect 10977 9129 11011 9163
rect 3157 9061 3191 9095
rect 10793 9061 10827 9095
rect 8493 8993 8527 9027
rect 16497 8993 16531 9027
rect 1593 8925 1627 8959
rect 1869 8925 1903 8959
rect 1961 8925 1995 8959
rect 2881 8925 2915 8959
rect 2973 8925 3007 8959
rect 3249 8925 3283 8959
rect 3341 8925 3375 8959
rect 4445 8925 4479 8959
rect 4813 8925 4847 8959
rect 4905 8925 4939 8959
rect 5089 8925 5123 8959
rect 5181 8925 5215 8959
rect 7573 8925 7607 8959
rect 16589 8925 16623 8959
rect 16960 8925 16994 8959
rect 17509 8925 17543 8959
rect 17693 8925 17727 8959
rect 18245 8925 18279 8959
rect 2237 8857 2271 8891
rect 3525 8857 3559 8891
rect 3893 8857 3927 8891
rect 8953 8857 8987 8891
rect 10945 8857 10979 8891
rect 11161 8857 11195 8891
rect 1777 8789 1811 8823
rect 5365 8789 5399 8823
rect 10425 8789 10459 8823
rect 16957 8789 16991 8823
rect 17141 8789 17175 8823
rect 17601 8789 17635 8823
rect 18429 8789 18463 8823
rect 2145 8585 2179 8619
rect 2329 8585 2363 8619
rect 7021 8585 7055 8619
rect 9413 8585 9447 8619
rect 10057 8585 10091 8619
rect 10425 8585 10459 8619
rect 1961 8517 1995 8551
rect 4537 8517 4571 8551
rect 10609 8517 10643 8551
rect 2237 8449 2271 8483
rect 3065 8449 3099 8483
rect 3157 8449 3191 8483
rect 4813 8449 4847 8483
rect 4997 8449 5031 8483
rect 5365 8449 5399 8483
rect 5549 8449 5583 8483
rect 6377 8449 6411 8483
rect 6561 8449 6595 8483
rect 6653 8449 6687 8483
rect 6745 8449 6779 8483
rect 7205 8449 7239 8483
rect 7389 8449 7423 8483
rect 9321 8449 9355 8483
rect 10149 8449 10183 8483
rect 10333 8449 10367 8483
rect 16681 8449 16715 8483
rect 16957 8449 16991 8483
rect 17049 8449 17083 8483
rect 2605 8381 2639 8415
rect 3746 8381 3780 8415
rect 6009 8381 6043 8415
rect 2513 8313 2547 8347
rect 6929 8313 6963 8347
rect 10609 8313 10643 8347
rect 3341 8245 3375 8279
rect 16773 8245 16807 8279
rect 17233 8245 17267 8279
rect 6009 8041 6043 8075
rect 13115 8041 13149 8075
rect 15761 8041 15795 8075
rect 1685 7973 1719 8007
rect 2513 7973 2547 8007
rect 13277 7973 13311 8007
rect 7205 7905 7239 7939
rect 9689 7905 9723 7939
rect 1409 7837 1443 7871
rect 4537 7837 4571 7871
rect 5825 7837 5859 7871
rect 6009 7837 6043 7871
rect 6561 7837 6595 7871
rect 6745 7837 6779 7871
rect 6837 7837 6871 7871
rect 6929 7837 6963 7871
rect 9229 7837 9263 7871
rect 9321 7837 9355 7871
rect 9597 7837 9631 7871
rect 9781 7837 9815 7871
rect 15117 7837 15151 7871
rect 15209 7837 15243 7871
rect 15393 7837 15427 7871
rect 15485 7837 15519 7871
rect 15577 7837 15611 7871
rect 15853 7837 15887 7871
rect 15945 7837 15979 7871
rect 16129 7837 16163 7871
rect 17509 7837 17543 7871
rect 18061 7837 18095 7871
rect 2697 7769 2731 7803
rect 2881 7769 2915 7803
rect 4353 7769 4387 7803
rect 9505 7769 9539 7803
rect 12909 7769 12943 7803
rect 13125 7769 13159 7803
rect 17325 7769 17359 7803
rect 1869 7701 1903 7735
rect 16313 7701 16347 7735
rect 9413 7497 9447 7531
rect 8217 7429 8251 7463
rect 7481 7361 7515 7395
rect 7573 7361 7607 7395
rect 7757 7361 7791 7395
rect 8769 7361 8803 7395
rect 9045 7361 9079 7395
rect 9873 7361 9907 7395
rect 10149 7361 10183 7395
rect 10333 7361 10367 7395
rect 10885 7361 10919 7395
rect 11529 7361 11563 7395
rect 11713 7361 11747 7395
rect 14197 7361 14231 7395
rect 14381 7361 14415 7395
rect 14657 7361 14691 7395
rect 17049 7361 17083 7395
rect 4261 7293 4295 7327
rect 4537 7293 4571 7327
rect 9965 7293 9999 7327
rect 11897 7293 11931 7327
rect 11069 7157 11103 7191
rect 17141 7157 17175 7191
rect 7849 6953 7883 6987
rect 12909 6885 12943 6919
rect 1685 6817 1719 6851
rect 4537 6817 4571 6851
rect 5089 6817 5123 6851
rect 3893 6749 3927 6783
rect 4077 6749 4111 6783
rect 4445 6749 4479 6783
rect 6653 6749 6687 6783
rect 7665 6749 7699 6783
rect 8033 6749 8067 6783
rect 8125 6749 8159 6783
rect 8217 6749 8251 6783
rect 8401 6749 8435 6783
rect 12633 6749 12667 6783
rect 18245 6749 18279 6783
rect 1501 6681 1535 6715
rect 13093 6613 13127 6647
rect 18429 6613 18463 6647
rect 4245 6409 4279 6443
rect 8217 6409 8251 6443
rect 9781 6409 9815 6443
rect 12357 6409 12391 6443
rect 3433 6341 3467 6375
rect 4445 6341 4479 6375
rect 7849 6341 7883 6375
rect 9873 6341 9907 6375
rect 10241 6341 10275 6375
rect 3617 6273 3651 6307
rect 3709 6273 3743 6307
rect 3893 6273 3927 6307
rect 3985 6273 4019 6307
rect 4813 6273 4847 6307
rect 4997 6273 5031 6307
rect 5273 6273 5307 6307
rect 5549 6273 5583 6307
rect 5733 6273 5767 6307
rect 8033 6273 8067 6307
rect 8125 6273 8159 6307
rect 9689 6273 9723 6307
rect 12173 6273 12207 6307
rect 12357 6273 12391 6307
rect 8401 6205 8435 6239
rect 9505 6205 9539 6239
rect 4077 6137 4111 6171
rect 4261 6069 4295 6103
rect 4905 6069 4939 6103
rect 5641 6069 5675 6103
rect 2605 5865 2639 5899
rect 6285 5865 6319 5899
rect 8953 5865 8987 5899
rect 10517 5865 10551 5899
rect 12449 5865 12483 5899
rect 17233 5865 17267 5899
rect 18061 5865 18095 5899
rect 7481 5797 7515 5831
rect 11069 5797 11103 5831
rect 2697 5729 2731 5763
rect 3065 5729 3099 5763
rect 3893 5729 3927 5763
rect 4353 5729 4387 5763
rect 6653 5729 6687 5763
rect 11621 5729 11655 5763
rect 14381 5729 14415 5763
rect 14473 5729 14507 5763
rect 14841 5729 14875 5763
rect 16589 5729 16623 5763
rect 2421 5661 2455 5695
rect 2513 5661 2547 5695
rect 4169 5661 4203 5695
rect 6561 5661 6595 5695
rect 7481 5661 7515 5695
rect 7757 5661 7791 5695
rect 9137 5661 9171 5695
rect 9505 5661 9539 5695
rect 10517 5661 10551 5695
rect 10793 5661 10827 5695
rect 11253 5661 11287 5695
rect 11345 5661 11379 5695
rect 11805 5661 11839 5695
rect 12541 5661 12575 5695
rect 14565 5661 14599 5695
rect 14657 5661 14691 5695
rect 15209 5661 15243 5695
rect 15577 5661 15611 5695
rect 16681 5661 16715 5695
rect 16773 5661 16807 5695
rect 16865 5661 16899 5695
rect 17601 5661 17635 5695
rect 17877 5661 17911 5695
rect 3801 5593 3835 5627
rect 9229 5593 9263 5627
rect 9321 5593 9355 5627
rect 10701 5593 10735 5627
rect 17693 5593 17727 5627
rect 3525 5525 3559 5559
rect 11437 5525 11471 5559
rect 14197 5525 14231 5559
rect 16405 5525 16439 5559
rect 7297 5321 7331 5355
rect 17509 5321 17543 5355
rect 8861 5253 8895 5287
rect 12633 5253 12667 5287
rect 16681 5253 16715 5287
rect 16865 5253 16899 5287
rect 3157 5185 3191 5219
rect 3801 5185 3835 5219
rect 4169 5185 4203 5219
rect 4445 5185 4479 5219
rect 4710 5185 4744 5219
rect 4997 5185 5031 5219
rect 5181 5185 5215 5219
rect 5641 5185 5675 5219
rect 6377 5185 6411 5219
rect 6561 5185 6595 5219
rect 6929 5185 6963 5219
rect 7665 5185 7699 5219
rect 7941 5185 7975 5219
rect 8309 5185 8343 5219
rect 9045 5185 9079 5219
rect 11897 5185 11931 5219
rect 12357 5185 12391 5219
rect 12449 5185 12483 5219
rect 15485 5185 15519 5219
rect 15669 5185 15703 5219
rect 17417 5185 17451 5219
rect 17601 5185 17635 5219
rect 18337 5185 18371 5219
rect 18521 5185 18555 5219
rect 4077 5117 4111 5151
rect 7021 5117 7055 5151
rect 7849 5117 7883 5151
rect 9229 5117 9263 5151
rect 11713 5117 11747 5151
rect 12081 5117 12115 5151
rect 16497 5117 16531 5151
rect 4813 5049 4847 5083
rect 5733 4981 5767 5015
rect 6101 4981 6135 5015
rect 12633 4981 12667 5015
rect 17049 4981 17083 5015
rect 18337 4981 18371 5015
rect 5273 4777 5307 4811
rect 5733 4777 5767 4811
rect 7849 4777 7883 4811
rect 11989 4777 12023 4811
rect 14657 4777 14691 4811
rect 2789 4709 2823 4743
rect 5365 4709 5399 4743
rect 7573 4709 7607 4743
rect 14473 4709 14507 4743
rect 3893 4641 3927 4675
rect 4353 4641 4387 4675
rect 4905 4641 4939 4675
rect 5089 4641 5123 4675
rect 7113 4641 7147 4675
rect 15577 4641 15611 4675
rect 1685 4573 1719 4607
rect 2053 4573 2087 4607
rect 2329 4573 2363 4607
rect 2881 4573 2915 4607
rect 3985 4573 4019 4607
rect 4813 4573 4847 4607
rect 4997 4573 5031 4607
rect 5549 4573 5583 4607
rect 5825 4573 5859 4607
rect 7205 4573 7239 4607
rect 7297 4573 7331 4607
rect 7389 4573 7423 4607
rect 7653 4573 7687 4607
rect 7849 4573 7883 4607
rect 10425 4573 10459 4607
rect 11253 4573 11287 4607
rect 11529 4573 11563 4607
rect 11805 4573 11839 4607
rect 14289 4573 14323 4607
rect 14565 4573 14599 4607
rect 14657 4573 14691 4607
rect 14841 4573 14875 4607
rect 15025 4573 15059 4607
rect 15209 4573 15243 4607
rect 14381 4505 14415 4539
rect 11621 4437 11655 4471
rect 2329 4233 2363 4267
rect 5641 4233 5675 4267
rect 5825 4165 5859 4199
rect 8493 4165 8527 4199
rect 16773 4165 16807 4199
rect 2053 4097 2087 4131
rect 2697 4097 2731 4131
rect 3341 4097 3375 4131
rect 3709 4097 3743 4131
rect 3985 4097 4019 4131
rect 4353 4097 4387 4131
rect 4629 4097 4663 4131
rect 5273 4097 5307 4131
rect 9137 4097 9171 4131
rect 9689 4097 9723 4131
rect 9873 4097 9907 4131
rect 12081 4097 12115 4131
rect 12173 4097 12207 4131
rect 12265 4097 12299 4131
rect 12449 4097 12483 4131
rect 12633 4097 12667 4131
rect 18245 4097 18279 4131
rect 1869 4029 1903 4063
rect 2421 4029 2455 4063
rect 2513 4029 2547 4063
rect 5181 4029 5215 4063
rect 9597 4029 9631 4063
rect 9781 4029 9815 4063
rect 10057 4029 10091 4063
rect 11989 4029 12023 4063
rect 12541 4029 12575 4063
rect 5457 3893 5491 3927
rect 5641 3893 5675 3927
rect 11805 3893 11839 3927
rect 16865 3893 16899 3927
rect 18429 3893 18463 3927
rect 6929 3689 6963 3723
rect 17141 3689 17175 3723
rect 17877 3689 17911 3723
rect 18061 3689 18095 3723
rect 8953 3621 8987 3655
rect 12909 3621 12943 3655
rect 1685 3553 1719 3587
rect 15945 3553 15979 3587
rect 17417 3553 17451 3587
rect 1409 3485 1443 3519
rect 2053 3485 2087 3519
rect 2697 3485 2731 3519
rect 2789 3485 2823 3519
rect 3065 3485 3099 3519
rect 4169 3485 4203 3519
rect 4353 3485 4387 3519
rect 4537 3485 4571 3519
rect 4629 3495 4663 3529
rect 6009 3485 6043 3519
rect 6193 3485 6227 3519
rect 7061 3485 7095 3519
rect 7205 3485 7239 3519
rect 7481 3485 7515 3519
rect 7941 3485 7975 3519
rect 8217 3485 8251 3519
rect 8309 3485 8343 3519
rect 8585 3485 8619 3519
rect 9137 3485 9171 3519
rect 9321 3485 9355 3519
rect 9413 3485 9447 3519
rect 12633 3485 12667 3519
rect 12725 3485 12759 3519
rect 13001 3485 13035 3519
rect 16037 3485 16071 3519
rect 16405 3485 16439 3519
rect 16497 3485 16531 3519
rect 16681 3485 16715 3519
rect 16865 3485 16899 3519
rect 17049 3485 17083 3519
rect 17233 3485 17267 3519
rect 17325 3485 17359 3519
rect 17601 3485 17635 3519
rect 17693 3485 17727 3519
rect 17969 3485 18003 3519
rect 18153 3485 18187 3519
rect 4261 3417 4295 3451
rect 6377 3417 6411 3451
rect 7297 3417 7331 3451
rect 8769 3417 8803 3451
rect 15393 3417 15427 3451
rect 2513 3349 2547 3383
rect 3985 3349 4019 3383
rect 7757 3349 7791 3383
rect 8125 3349 8159 3383
rect 8401 3349 8435 3383
rect 12449 3349 12483 3383
rect 16773 3349 16807 3383
rect 3433 3145 3467 3179
rect 8953 3145 8987 3179
rect 11697 3145 11731 3179
rect 1777 3077 1811 3111
rect 5365 3077 5399 3111
rect 11345 3077 11379 3111
rect 11897 3077 11931 3111
rect 12173 3077 12207 3111
rect 2421 3009 2455 3043
rect 2789 3009 2823 3043
rect 2973 3009 3007 3043
rect 3065 3009 3099 3043
rect 3525 3009 3559 3043
rect 6377 3009 6411 3043
rect 6561 3009 6595 3043
rect 6837 3009 6871 3043
rect 8125 3009 8159 3043
rect 8309 3009 8343 3043
rect 8401 3031 8435 3065
rect 8493 3009 8527 3043
rect 8769 3009 8803 3043
rect 9321 3009 9355 3043
rect 9413 3009 9447 3043
rect 9597 3009 9631 3043
rect 9781 3009 9815 3043
rect 11161 3009 11195 3043
rect 12081 3009 12115 3043
rect 12265 3009 12299 3043
rect 13093 3009 13127 3043
rect 17233 3009 17267 3043
rect 17417 3009 17451 3043
rect 2237 2941 2271 2975
rect 3157 2941 3191 2975
rect 3249 2941 3283 2975
rect 7941 2941 7975 2975
rect 8585 2941 8619 2975
rect 12725 2941 12759 2975
rect 13277 2941 13311 2975
rect 1593 2873 1627 2907
rect 2697 2873 2731 2907
rect 3893 2873 3927 2907
rect 6653 2873 6687 2907
rect 6745 2873 6779 2907
rect 12817 2873 12851 2907
rect 3985 2805 4019 2839
rect 5273 2805 5307 2839
rect 7021 2805 7055 2839
rect 11069 2805 11103 2839
rect 11529 2805 11563 2839
rect 11713 2805 11747 2839
rect 17325 2805 17359 2839
rect 2329 2601 2363 2635
rect 2789 2601 2823 2635
rect 3985 2601 4019 2635
rect 6653 2601 6687 2635
rect 9045 2601 9079 2635
rect 12817 2533 12851 2567
rect 1409 2465 1443 2499
rect 2513 2465 2547 2499
rect 8125 2465 8159 2499
rect 8585 2465 8619 2499
rect 8677 2465 8711 2499
rect 9505 2465 9539 2499
rect 10425 2465 10459 2499
rect 12357 2465 12391 2499
rect 1869 2397 1903 2431
rect 1961 2397 1995 2431
rect 2053 2397 2087 2431
rect 2237 2397 2271 2431
rect 2605 2397 2639 2431
rect 6561 2397 6595 2431
rect 7080 2397 7114 2431
rect 8309 2397 8343 2431
rect 9229 2397 9263 2431
rect 9321 2397 9355 2431
rect 9597 2397 9631 2431
rect 11161 2397 11195 2431
rect 11345 2397 11379 2431
rect 11805 2397 11839 2431
rect 11989 2397 12023 2431
rect 12081 2397 12115 2431
rect 12633 2397 12667 2431
rect 12909 2397 12943 2431
rect 16681 2397 16715 2431
rect 17509 2397 17543 2431
rect 3893 2329 3927 2363
rect 10149 2329 10183 2363
rect 18337 2329 18371 2363
rect 2513 2261 2547 2295
rect 7021 2261 7055 2295
rect 7205 2261 7239 2295
rect 11161 2261 11195 2295
rect 11621 2261 11655 2295
rect 16865 2261 16899 2295
<< metal1 >>
rect 5810 18776 5816 18828
rect 5868 18816 5874 18828
rect 11514 18816 11520 18828
rect 5868 18788 11520 18816
rect 5868 18776 5874 18788
rect 11514 18776 11520 18788
rect 11572 18776 11578 18828
rect 6086 18708 6092 18760
rect 6144 18748 6150 18760
rect 14274 18748 14280 18760
rect 6144 18720 14280 18748
rect 6144 18708 6150 18720
rect 14274 18708 14280 18720
rect 14332 18708 14338 18760
rect 1578 18572 1584 18624
rect 1636 18612 1642 18624
rect 10226 18612 10232 18624
rect 1636 18584 10232 18612
rect 1636 18572 1642 18584
rect 10226 18572 10232 18584
rect 10284 18572 10290 18624
rect 5626 18504 5632 18556
rect 5684 18544 5690 18556
rect 15930 18544 15936 18556
rect 5684 18516 15936 18544
rect 5684 18504 5690 18516
rect 15930 18504 15936 18516
rect 15988 18504 15994 18556
rect 3326 18436 3332 18488
rect 3384 18476 3390 18488
rect 14458 18476 14464 18488
rect 3384 18448 14464 18476
rect 3384 18436 3390 18448
rect 14458 18436 14464 18448
rect 14516 18436 14522 18488
rect 9674 18368 9680 18420
rect 9732 18408 9738 18420
rect 11422 18408 11428 18420
rect 9732 18380 11428 18408
rect 9732 18368 9738 18380
rect 11422 18368 11428 18380
rect 11480 18368 11486 18420
rect 11514 18368 11520 18420
rect 11572 18408 11578 18420
rect 16758 18408 16764 18420
rect 11572 18380 16764 18408
rect 11572 18368 11578 18380
rect 16758 18368 16764 18380
rect 16816 18368 16822 18420
rect 5258 18300 5264 18352
rect 5316 18340 5322 18352
rect 14642 18340 14648 18352
rect 5316 18312 14648 18340
rect 5316 18300 5322 18312
rect 14642 18300 14648 18312
rect 14700 18300 14706 18352
rect 8570 18232 8576 18284
rect 8628 18272 8634 18284
rect 14366 18272 14372 18284
rect 8628 18244 14372 18272
rect 8628 18232 8634 18244
rect 14366 18232 14372 18244
rect 14424 18232 14430 18284
rect 6730 18164 6736 18216
rect 6788 18204 6794 18216
rect 6788 18176 6914 18204
rect 6788 18164 6794 18176
rect 6886 18136 6914 18176
rect 11422 18164 11428 18216
rect 11480 18204 11486 18216
rect 16298 18204 16304 18216
rect 11480 18176 16304 18204
rect 11480 18164 11486 18176
rect 16298 18164 16304 18176
rect 16356 18164 16362 18216
rect 13814 18136 13820 18148
rect 6886 18108 13820 18136
rect 13814 18096 13820 18108
rect 13872 18096 13878 18148
rect 9030 18028 9036 18080
rect 9088 18068 9094 18080
rect 15286 18068 15292 18080
rect 9088 18040 15292 18068
rect 9088 18028 9094 18040
rect 15286 18028 15292 18040
rect 15344 18028 15350 18080
rect 3602 17960 3608 18012
rect 3660 18000 3666 18012
rect 10778 18000 10784 18012
rect 3660 17972 10784 18000
rect 3660 17960 3666 17972
rect 10778 17960 10784 17972
rect 10836 17960 10842 18012
rect 4430 17756 4436 17808
rect 4488 17796 4494 17808
rect 9582 17796 9588 17808
rect 4488 17768 9588 17796
rect 4488 17756 4494 17768
rect 9582 17756 9588 17768
rect 9640 17756 9646 17808
rect 15930 17756 15936 17808
rect 15988 17796 15994 17808
rect 19518 17796 19524 17808
rect 15988 17768 19524 17796
rect 15988 17756 15994 17768
rect 19518 17756 19524 17768
rect 19576 17756 19582 17808
rect 4798 17688 4804 17740
rect 4856 17728 4862 17740
rect 9858 17728 9864 17740
rect 4856 17700 9864 17728
rect 4856 17688 4862 17700
rect 9858 17688 9864 17700
rect 9916 17688 9922 17740
rect 3970 17620 3976 17672
rect 4028 17660 4034 17672
rect 16482 17660 16488 17672
rect 4028 17632 16488 17660
rect 4028 17620 4034 17632
rect 16482 17620 16488 17632
rect 16540 17620 16546 17672
rect 8202 17552 8208 17604
rect 8260 17592 8266 17604
rect 15378 17592 15384 17604
rect 8260 17564 15384 17592
rect 8260 17552 8266 17564
rect 15378 17552 15384 17564
rect 15436 17552 15442 17604
rect 3510 17484 3516 17536
rect 3568 17524 3574 17536
rect 9766 17524 9772 17536
rect 3568 17496 9772 17524
rect 3568 17484 3574 17496
rect 9766 17484 9772 17496
rect 9824 17484 9830 17536
rect 9858 17484 9864 17536
rect 9916 17524 9922 17536
rect 16666 17524 16672 17536
rect 9916 17496 16672 17524
rect 9916 17484 9922 17496
rect 16666 17484 16672 17496
rect 16724 17484 16730 17536
rect 1104 17434 18860 17456
rect 1104 17382 2610 17434
rect 2662 17382 2674 17434
rect 2726 17382 2738 17434
rect 2790 17382 2802 17434
rect 2854 17382 2866 17434
rect 2918 17382 7610 17434
rect 7662 17382 7674 17434
rect 7726 17382 7738 17434
rect 7790 17382 7802 17434
rect 7854 17382 7866 17434
rect 7918 17382 12610 17434
rect 12662 17382 12674 17434
rect 12726 17382 12738 17434
rect 12790 17382 12802 17434
rect 12854 17382 12866 17434
rect 12918 17382 17610 17434
rect 17662 17382 17674 17434
rect 17726 17382 17738 17434
rect 17790 17382 17802 17434
rect 17854 17382 17866 17434
rect 17918 17382 18860 17434
rect 1104 17360 18860 17382
rect 934 17280 940 17332
rect 992 17320 998 17332
rect 9033 17323 9091 17329
rect 9033 17320 9045 17323
rect 992 17292 9045 17320
rect 992 17280 998 17292
rect 9033 17289 9045 17292
rect 9079 17289 9091 17323
rect 9033 17283 9091 17289
rect 9490 17280 9496 17332
rect 9548 17320 9554 17332
rect 15654 17320 15660 17332
rect 9548 17292 15660 17320
rect 9548 17280 9554 17292
rect 15654 17280 15660 17292
rect 15712 17280 15718 17332
rect 17494 17280 17500 17332
rect 17552 17320 17558 17332
rect 17865 17323 17923 17329
rect 17865 17320 17877 17323
rect 17552 17292 17877 17320
rect 17552 17280 17558 17292
rect 17865 17289 17877 17292
rect 17911 17289 17923 17323
rect 17865 17283 17923 17289
rect 2409 17255 2467 17261
rect 2409 17221 2421 17255
rect 2455 17252 2467 17255
rect 2958 17252 2964 17264
rect 2455 17224 2964 17252
rect 2455 17221 2467 17224
rect 2409 17215 2467 17221
rect 2958 17212 2964 17224
rect 3016 17212 3022 17264
rect 3694 17212 3700 17264
rect 3752 17252 3758 17264
rect 3881 17255 3939 17261
rect 3881 17252 3893 17255
rect 3752 17224 3893 17252
rect 3752 17212 3758 17224
rect 3881 17221 3893 17224
rect 3927 17221 3939 17255
rect 3881 17215 3939 17221
rect 4249 17255 4307 17261
rect 4249 17221 4261 17255
rect 4295 17252 4307 17255
rect 4295 17224 6132 17252
rect 4295 17221 4307 17224
rect 4249 17215 4307 17221
rect 2225 17187 2283 17193
rect 2225 17153 2237 17187
rect 2271 17184 2283 17187
rect 3050 17184 3056 17196
rect 2271 17156 3056 17184
rect 2271 17153 2283 17156
rect 2225 17147 2283 17153
rect 3050 17144 3056 17156
rect 3108 17144 3114 17196
rect 5442 17144 5448 17196
rect 5500 17144 5506 17196
rect 6104 17184 6132 17224
rect 6178 17212 6184 17264
rect 6236 17252 6242 17264
rect 6457 17255 6515 17261
rect 6457 17252 6469 17255
rect 6236 17224 6469 17252
rect 6236 17212 6242 17224
rect 6457 17221 6469 17224
rect 6503 17221 6515 17255
rect 6457 17215 6515 17221
rect 8662 17212 8668 17264
rect 8720 17252 8726 17264
rect 9585 17255 9643 17261
rect 9585 17252 9597 17255
rect 8720 17224 9597 17252
rect 8720 17212 8726 17224
rect 9585 17221 9597 17224
rect 9631 17221 9643 17255
rect 9585 17215 9643 17221
rect 9766 17212 9772 17264
rect 9824 17212 9830 17264
rect 13170 17252 13176 17264
rect 10888 17224 13176 17252
rect 7374 17184 7380 17196
rect 6104 17156 7380 17184
rect 7374 17144 7380 17156
rect 7432 17144 7438 17196
rect 9217 17187 9275 17193
rect 9217 17153 9229 17187
rect 9263 17153 9275 17187
rect 9217 17147 9275 17153
rect 9401 17187 9459 17193
rect 9401 17153 9413 17187
rect 9447 17184 9459 17187
rect 10888 17184 10916 17224
rect 13170 17212 13176 17224
rect 13228 17212 13234 17264
rect 9447 17156 10916 17184
rect 11057 17187 11115 17193
rect 9447 17153 9459 17156
rect 9401 17147 9459 17153
rect 11057 17153 11069 17187
rect 11103 17184 11115 17187
rect 11146 17184 11152 17196
rect 11103 17156 11152 17184
rect 11103 17153 11115 17156
rect 11057 17147 11115 17153
rect 5350 17076 5356 17128
rect 5408 17076 5414 17128
rect 9232 17116 9260 17147
rect 11146 17144 11152 17156
rect 11204 17144 11210 17196
rect 11793 17187 11851 17193
rect 11793 17153 11805 17187
rect 11839 17153 11851 17187
rect 11793 17147 11851 17153
rect 9582 17116 9588 17128
rect 9232 17088 9588 17116
rect 9582 17076 9588 17088
rect 9640 17076 9646 17128
rect 10502 17076 10508 17128
rect 10560 17116 10566 17128
rect 11808 17116 11836 17147
rect 13630 17144 13636 17196
rect 13688 17184 13694 17196
rect 14093 17187 14151 17193
rect 14093 17184 14105 17187
rect 13688 17156 14105 17184
rect 13688 17144 13694 17156
rect 14093 17153 14105 17156
rect 14139 17153 14151 17187
rect 14093 17147 14151 17153
rect 16114 17144 16120 17196
rect 16172 17184 16178 17196
rect 16393 17187 16451 17193
rect 16393 17184 16405 17187
rect 16172 17156 16405 17184
rect 16172 17144 16178 17156
rect 16393 17153 16405 17156
rect 16439 17153 16451 17187
rect 16393 17147 16451 17153
rect 17310 17144 17316 17196
rect 17368 17184 17374 17196
rect 17681 17187 17739 17193
rect 17681 17184 17693 17187
rect 17368 17156 17693 17184
rect 17368 17144 17374 17156
rect 17681 17153 17693 17156
rect 17727 17153 17739 17187
rect 17681 17147 17739 17153
rect 18509 17187 18567 17193
rect 18509 17153 18521 17187
rect 18555 17184 18567 17187
rect 18598 17184 18604 17196
rect 18555 17156 18604 17184
rect 18555 17153 18567 17156
rect 18509 17147 18567 17153
rect 18598 17144 18604 17156
rect 18656 17144 18662 17196
rect 10560 17088 11836 17116
rect 11885 17119 11943 17125
rect 10560 17076 10566 17088
rect 11885 17085 11897 17119
rect 11931 17085 11943 17119
rect 11885 17079 11943 17085
rect 5813 17051 5871 17057
rect 5813 17017 5825 17051
rect 5859 17048 5871 17051
rect 10410 17048 10416 17060
rect 5859 17020 10416 17048
rect 5859 17017 5871 17020
rect 5813 17011 5871 17017
rect 10410 17008 10416 17020
rect 10468 17008 10474 17060
rect 11900 17048 11928 17079
rect 11974 17076 11980 17128
rect 12032 17116 12038 17128
rect 12621 17119 12679 17125
rect 12621 17116 12633 17119
rect 12032 17088 12633 17116
rect 12032 17076 12038 17088
rect 12621 17085 12633 17088
rect 12667 17085 12679 17119
rect 12621 17079 12679 17085
rect 10888 17020 11928 17048
rect 12636 17048 12664 17079
rect 16022 17076 16028 17128
rect 16080 17076 16086 17128
rect 18138 17076 18144 17128
rect 18196 17116 18202 17128
rect 18233 17119 18291 17125
rect 18233 17116 18245 17119
rect 18196 17088 18245 17116
rect 18196 17076 18202 17088
rect 18233 17085 18245 17088
rect 18279 17085 18291 17119
rect 18233 17079 18291 17085
rect 17310 17048 17316 17060
rect 12636 17020 17316 17048
rect 1762 16940 1768 16992
rect 1820 16940 1826 16992
rect 2133 16983 2191 16989
rect 2133 16949 2145 16983
rect 2179 16980 2191 16983
rect 2406 16980 2412 16992
rect 2179 16952 2412 16980
rect 2179 16949 2191 16952
rect 2133 16943 2191 16949
rect 2406 16940 2412 16952
rect 2464 16980 2470 16992
rect 2501 16983 2559 16989
rect 2501 16980 2513 16983
rect 2464 16952 2513 16980
rect 2464 16940 2470 16952
rect 2501 16949 2513 16952
rect 2547 16949 2559 16983
rect 2501 16943 2559 16949
rect 4890 16940 4896 16992
rect 4948 16980 4954 16992
rect 6270 16980 6276 16992
rect 4948 16952 6276 16980
rect 4948 16940 4954 16952
rect 6270 16940 6276 16952
rect 6328 16980 6334 16992
rect 6549 16983 6607 16989
rect 6549 16980 6561 16983
rect 6328 16952 6561 16980
rect 6328 16940 6334 16952
rect 6549 16949 6561 16952
rect 6595 16949 6607 16983
rect 6549 16943 6607 16949
rect 8754 16940 8760 16992
rect 8812 16980 8818 16992
rect 10888 16980 10916 17020
rect 17310 17008 17316 17020
rect 17368 17008 17374 17060
rect 8812 16952 10916 16980
rect 11241 16983 11299 16989
rect 8812 16940 8818 16952
rect 11241 16949 11253 16983
rect 11287 16980 11299 16983
rect 11330 16980 11336 16992
rect 11287 16952 11336 16980
rect 11287 16949 11299 16952
rect 11241 16943 11299 16949
rect 11330 16940 11336 16952
rect 11388 16940 11394 16992
rect 12986 16940 12992 16992
rect 13044 16980 13050 16992
rect 14277 16983 14335 16989
rect 14277 16980 14289 16983
rect 13044 16952 14289 16980
rect 13044 16940 13050 16952
rect 14277 16949 14289 16952
rect 14323 16949 14335 16983
rect 14277 16943 14335 16949
rect 1104 16890 18860 16912
rect 1104 16838 1950 16890
rect 2002 16838 2014 16890
rect 2066 16838 2078 16890
rect 2130 16838 2142 16890
rect 2194 16838 2206 16890
rect 2258 16838 6950 16890
rect 7002 16838 7014 16890
rect 7066 16838 7078 16890
rect 7130 16838 7142 16890
rect 7194 16838 7206 16890
rect 7258 16838 11950 16890
rect 12002 16838 12014 16890
rect 12066 16838 12078 16890
rect 12130 16838 12142 16890
rect 12194 16838 12206 16890
rect 12258 16838 16950 16890
rect 17002 16838 17014 16890
rect 17066 16838 17078 16890
rect 17130 16838 17142 16890
rect 17194 16838 17206 16890
rect 17258 16838 18860 16890
rect 1104 16816 18860 16838
rect 8110 16736 8116 16788
rect 8168 16776 8174 16788
rect 13538 16776 13544 16788
rect 8168 16748 13544 16776
rect 8168 16736 8174 16748
rect 13538 16736 13544 16748
rect 13596 16736 13602 16788
rect 13722 16736 13728 16788
rect 13780 16776 13786 16788
rect 13780 16748 15332 16776
rect 13780 16736 13786 16748
rect 4982 16668 4988 16720
rect 5040 16708 5046 16720
rect 10502 16708 10508 16720
rect 5040 16680 10508 16708
rect 5040 16668 5046 16680
rect 10502 16668 10508 16680
rect 10560 16668 10566 16720
rect 10686 16668 10692 16720
rect 10744 16668 10750 16720
rect 10778 16668 10784 16720
rect 10836 16708 10842 16720
rect 14829 16711 14887 16717
rect 14829 16708 14841 16711
rect 10836 16680 14841 16708
rect 10836 16668 10842 16680
rect 14829 16677 14841 16680
rect 14875 16677 14887 16711
rect 14829 16671 14887 16677
rect 1854 16600 1860 16652
rect 1912 16640 1918 16652
rect 2225 16643 2283 16649
rect 2225 16640 2237 16643
rect 1912 16612 2237 16640
rect 1912 16600 1918 16612
rect 2225 16609 2237 16612
rect 2271 16609 2283 16643
rect 2225 16603 2283 16609
rect 5442 16600 5448 16652
rect 5500 16640 5506 16652
rect 8570 16640 8576 16652
rect 5500 16612 8576 16640
rect 5500 16600 5506 16612
rect 8570 16600 8576 16612
rect 8628 16600 8634 16652
rect 8846 16600 8852 16652
rect 8904 16640 8910 16652
rect 10965 16643 11023 16649
rect 10965 16640 10977 16643
rect 8904 16612 10977 16640
rect 8904 16600 8910 16612
rect 10965 16609 10977 16612
rect 11011 16609 11023 16643
rect 10965 16603 11023 16609
rect 11333 16643 11391 16649
rect 11333 16609 11345 16643
rect 11379 16640 11391 16643
rect 12434 16640 12440 16652
rect 11379 16612 12440 16640
rect 11379 16609 11391 16612
rect 11333 16603 11391 16609
rect 12434 16600 12440 16612
rect 12492 16600 12498 16652
rect 15194 16600 15200 16652
rect 15252 16600 15258 16652
rect 15304 16640 15332 16748
rect 15562 16736 15568 16788
rect 15620 16776 15626 16788
rect 16577 16779 16635 16785
rect 16577 16776 16589 16779
rect 15620 16748 16589 16776
rect 15620 16736 15626 16748
rect 16577 16745 16589 16748
rect 16623 16745 16635 16779
rect 16577 16739 16635 16745
rect 16206 16668 16212 16720
rect 16264 16708 16270 16720
rect 16761 16711 16819 16717
rect 16761 16708 16773 16711
rect 16264 16680 16773 16708
rect 16264 16668 16270 16680
rect 16761 16677 16773 16680
rect 16807 16677 16819 16711
rect 16761 16671 16819 16677
rect 16853 16711 16911 16717
rect 16853 16677 16865 16711
rect 16899 16677 16911 16711
rect 16853 16671 16911 16677
rect 16868 16640 16896 16671
rect 15304 16612 16896 16640
rect 1210 16532 1216 16584
rect 1268 16572 1274 16584
rect 2041 16575 2099 16581
rect 2041 16572 2053 16575
rect 1268 16544 2053 16572
rect 1268 16532 1274 16544
rect 2041 16541 2053 16544
rect 2087 16541 2099 16575
rect 2041 16535 2099 16541
rect 10410 16532 10416 16584
rect 10468 16532 10474 16584
rect 10594 16532 10600 16584
rect 10652 16572 10658 16584
rect 11149 16575 11207 16581
rect 11149 16572 11161 16575
rect 10652 16544 11161 16572
rect 10652 16532 10658 16544
rect 11149 16541 11161 16544
rect 11195 16541 11207 16575
rect 11149 16535 11207 16541
rect 11606 16532 11612 16584
rect 11664 16572 11670 16584
rect 15105 16575 15163 16581
rect 15105 16572 15117 16575
rect 11664 16544 15117 16572
rect 11664 16532 11670 16544
rect 15105 16541 15117 16544
rect 15151 16541 15163 16575
rect 15105 16535 15163 16541
rect 16114 16532 16120 16584
rect 16172 16572 16178 16584
rect 16853 16575 16911 16581
rect 16853 16572 16865 16575
rect 16172 16544 16865 16572
rect 16172 16532 16178 16544
rect 16853 16541 16865 16544
rect 16899 16541 16911 16575
rect 16853 16535 16911 16541
rect 17034 16532 17040 16584
rect 17092 16532 17098 16584
rect 17126 16532 17132 16584
rect 17184 16532 17190 16584
rect 18233 16575 18291 16581
rect 18233 16541 18245 16575
rect 18279 16541 18291 16575
rect 18233 16535 18291 16541
rect 1486 16464 1492 16516
rect 1544 16464 1550 16516
rect 1857 16507 1915 16513
rect 1857 16473 1869 16507
rect 1903 16504 1915 16507
rect 3142 16504 3148 16516
rect 1903 16476 3148 16504
rect 1903 16473 1915 16476
rect 1857 16467 1915 16473
rect 3142 16464 3148 16476
rect 3200 16464 3206 16516
rect 10689 16507 10747 16513
rect 10689 16473 10701 16507
rect 10735 16504 10747 16507
rect 11330 16504 11336 16516
rect 10735 16476 11336 16504
rect 10735 16473 10747 16476
rect 10689 16467 10747 16473
rect 11330 16464 11336 16476
rect 11388 16464 11394 16516
rect 11514 16464 11520 16516
rect 11572 16504 11578 16516
rect 13446 16504 13452 16516
rect 11572 16476 13452 16504
rect 11572 16464 11578 16476
rect 13446 16464 13452 16476
rect 13504 16464 13510 16516
rect 14182 16464 14188 16516
rect 14240 16504 14246 16516
rect 14553 16507 14611 16513
rect 14553 16504 14565 16507
rect 14240 16476 14565 16504
rect 14240 16464 14246 16476
rect 14553 16473 14565 16476
rect 14599 16473 14611 16507
rect 14553 16467 14611 16473
rect 16390 16464 16396 16516
rect 16448 16464 16454 16516
rect 17954 16504 17960 16516
rect 16608 16476 17960 16504
rect 10502 16396 10508 16448
rect 10560 16396 10566 16448
rect 10870 16396 10876 16448
rect 10928 16436 10934 16448
rect 16608 16445 16636 16476
rect 17954 16464 17960 16476
rect 18012 16464 18018 16516
rect 16593 16439 16651 16445
rect 16593 16436 16605 16439
rect 10928 16408 16605 16436
rect 10928 16396 10934 16408
rect 16593 16405 16605 16408
rect 16639 16405 16651 16439
rect 16593 16399 16651 16405
rect 16758 16396 16764 16448
rect 16816 16436 16822 16448
rect 17865 16439 17923 16445
rect 17865 16436 17877 16439
rect 16816 16408 17877 16436
rect 16816 16396 16822 16408
rect 17865 16405 17877 16408
rect 17911 16436 17923 16439
rect 18248 16436 18276 16535
rect 17911 16408 18276 16436
rect 17911 16405 17923 16408
rect 17865 16399 17923 16405
rect 18414 16396 18420 16448
rect 18472 16396 18478 16448
rect 1104 16346 18860 16368
rect 1104 16294 2610 16346
rect 2662 16294 2674 16346
rect 2726 16294 2738 16346
rect 2790 16294 2802 16346
rect 2854 16294 2866 16346
rect 2918 16294 7610 16346
rect 7662 16294 7674 16346
rect 7726 16294 7738 16346
rect 7790 16294 7802 16346
rect 7854 16294 7866 16346
rect 7918 16294 12610 16346
rect 12662 16294 12674 16346
rect 12726 16294 12738 16346
rect 12790 16294 12802 16346
rect 12854 16294 12866 16346
rect 12918 16294 17610 16346
rect 17662 16294 17674 16346
rect 17726 16294 17738 16346
rect 17790 16294 17802 16346
rect 17854 16294 17866 16346
rect 17918 16294 18860 16346
rect 1104 16272 18860 16294
rect 3053 16235 3111 16241
rect 3053 16201 3065 16235
rect 3099 16232 3111 16235
rect 4614 16232 4620 16244
rect 3099 16204 4620 16232
rect 3099 16201 3111 16204
rect 3053 16195 3111 16201
rect 3068 16164 3096 16195
rect 4614 16192 4620 16204
rect 4672 16192 4678 16244
rect 5166 16192 5172 16244
rect 5224 16232 5230 16244
rect 12986 16232 12992 16244
rect 5224 16204 12992 16232
rect 5224 16192 5230 16204
rect 12986 16192 12992 16204
rect 13044 16192 13050 16244
rect 16945 16235 17003 16241
rect 16945 16201 16957 16235
rect 16991 16232 17003 16235
rect 17126 16232 17132 16244
rect 16991 16204 17132 16232
rect 16991 16201 17003 16204
rect 16945 16195 17003 16201
rect 17126 16192 17132 16204
rect 17184 16192 17190 16244
rect 2976 16136 3096 16164
rect 2685 16031 2743 16037
rect 2685 15997 2697 16031
rect 2731 16028 2743 16031
rect 2774 16028 2780 16040
rect 2731 16000 2780 16028
rect 2731 15997 2743 16000
rect 2685 15991 2743 15997
rect 2774 15988 2780 16000
rect 2832 15988 2838 16040
rect 842 15920 848 15972
rect 900 15960 906 15972
rect 2976 15960 3004 16136
rect 7374 16124 7380 16176
rect 7432 16164 7438 16176
rect 9122 16164 9128 16176
rect 7432 16136 9128 16164
rect 7432 16124 7438 16136
rect 9122 16124 9128 16136
rect 9180 16164 9186 16176
rect 9180 16136 12480 16164
rect 9180 16124 9186 16136
rect 3050 16056 3056 16108
rect 3108 16056 3114 16108
rect 6546 16056 6552 16108
rect 6604 16056 6610 16108
rect 6638 16056 6644 16108
rect 6696 16056 6702 16108
rect 7006 16056 7012 16108
rect 7064 16056 7070 16108
rect 7834 16056 7840 16108
rect 7892 16096 7898 16108
rect 8202 16096 8208 16108
rect 7892 16068 8208 16096
rect 7892 16056 7898 16068
rect 8202 16056 8208 16068
rect 8260 16056 8266 16108
rect 9214 16056 9220 16108
rect 9272 16096 9278 16108
rect 12161 16099 12219 16105
rect 12161 16096 12173 16099
rect 9272 16068 12173 16096
rect 9272 16056 9278 16068
rect 12161 16065 12173 16068
rect 12207 16065 12219 16099
rect 12161 16059 12219 16065
rect 12345 16099 12403 16105
rect 12345 16065 12357 16099
rect 12391 16065 12403 16099
rect 12452 16096 12480 16136
rect 12526 16124 12532 16176
rect 12584 16164 12590 16176
rect 12713 16167 12771 16173
rect 12713 16164 12725 16167
rect 12584 16136 12725 16164
rect 12584 16124 12590 16136
rect 12713 16133 12725 16136
rect 12759 16133 12771 16167
rect 12713 16127 12771 16133
rect 13538 16124 13544 16176
rect 13596 16164 13602 16176
rect 18230 16164 18236 16176
rect 13596 16136 18236 16164
rect 13596 16124 13602 16136
rect 18230 16124 18236 16136
rect 18288 16124 18294 16176
rect 12618 16096 12624 16108
rect 12452 16068 12624 16096
rect 12345 16059 12403 16065
rect 3237 16031 3295 16037
rect 3237 15997 3249 16031
rect 3283 16028 3295 16031
rect 6454 16028 6460 16040
rect 3283 16000 6460 16028
rect 3283 15997 3295 16000
rect 3237 15991 3295 15997
rect 6454 15988 6460 16000
rect 6512 15988 6518 16040
rect 7742 15988 7748 16040
rect 7800 16028 7806 16040
rect 10410 16028 10416 16040
rect 7800 16000 10416 16028
rect 7800 15988 7806 16000
rect 10410 15988 10416 16000
rect 10468 15988 10474 16040
rect 10870 15988 10876 16040
rect 10928 16028 10934 16040
rect 11606 16028 11612 16040
rect 10928 16000 11612 16028
rect 10928 15988 10934 16000
rect 11606 15988 11612 16000
rect 11664 15988 11670 16040
rect 12360 16028 12388 16059
rect 12618 16056 12624 16068
rect 12676 16056 12682 16108
rect 12897 16099 12955 16105
rect 12897 16065 12909 16099
rect 12943 16096 12955 16099
rect 16574 16096 16580 16108
rect 12943 16068 16580 16096
rect 12943 16065 12955 16068
rect 12897 16059 12955 16065
rect 16574 16056 16580 16068
rect 16632 16056 16638 16108
rect 17494 16028 17500 16040
rect 12360 16000 17500 16028
rect 17494 15988 17500 16000
rect 17552 15988 17558 16040
rect 900 15932 3004 15960
rect 900 15920 906 15932
rect 4154 15920 4160 15972
rect 4212 15960 4218 15972
rect 10042 15960 10048 15972
rect 4212 15932 10048 15960
rect 4212 15920 4218 15932
rect 10042 15920 10048 15932
rect 10100 15920 10106 15972
rect 10686 15920 10692 15972
rect 10744 15960 10750 15972
rect 12526 15960 12532 15972
rect 10744 15932 12532 15960
rect 10744 15920 10750 15932
rect 12526 15920 12532 15932
rect 12584 15920 12590 15972
rect 6917 15895 6975 15901
rect 6917 15861 6929 15895
rect 6963 15892 6975 15895
rect 7374 15892 7380 15904
rect 6963 15864 7380 15892
rect 6963 15861 6975 15864
rect 6917 15855 6975 15861
rect 7374 15852 7380 15864
rect 7432 15852 7438 15904
rect 8018 15852 8024 15904
rect 8076 15892 8082 15904
rect 10318 15892 10324 15904
rect 8076 15864 10324 15892
rect 8076 15852 8082 15864
rect 10318 15852 10324 15864
rect 10376 15852 10382 15904
rect 11606 15852 11612 15904
rect 11664 15892 11670 15904
rect 12253 15895 12311 15901
rect 12253 15892 12265 15895
rect 11664 15864 12265 15892
rect 11664 15852 11670 15864
rect 12253 15861 12265 15864
rect 12299 15861 12311 15895
rect 12253 15855 12311 15861
rect 12897 15895 12955 15901
rect 12897 15861 12909 15895
rect 12943 15892 12955 15895
rect 18782 15892 18788 15904
rect 12943 15864 18788 15892
rect 12943 15861 12955 15864
rect 12897 15855 12955 15861
rect 18782 15852 18788 15864
rect 18840 15852 18846 15904
rect 1104 15802 18860 15824
rect 1104 15750 1950 15802
rect 2002 15750 2014 15802
rect 2066 15750 2078 15802
rect 2130 15750 2142 15802
rect 2194 15750 2206 15802
rect 2258 15750 6950 15802
rect 7002 15750 7014 15802
rect 7066 15750 7078 15802
rect 7130 15750 7142 15802
rect 7194 15750 7206 15802
rect 7258 15750 11950 15802
rect 12002 15750 12014 15802
rect 12066 15750 12078 15802
rect 12130 15750 12142 15802
rect 12194 15750 12206 15802
rect 12258 15750 16950 15802
rect 17002 15750 17014 15802
rect 17066 15750 17078 15802
rect 17130 15750 17142 15802
rect 17194 15750 17206 15802
rect 17258 15750 18860 15802
rect 1104 15728 18860 15750
rect 1854 15648 1860 15700
rect 1912 15688 1918 15700
rect 5350 15688 5356 15700
rect 1912 15660 5356 15688
rect 1912 15648 1918 15660
rect 5350 15648 5356 15660
rect 5408 15648 5414 15700
rect 5442 15648 5448 15700
rect 5500 15648 5506 15700
rect 5718 15648 5724 15700
rect 5776 15688 5782 15700
rect 5776 15660 8340 15688
rect 5776 15648 5782 15660
rect 2774 15580 2780 15632
rect 2832 15620 2838 15632
rect 3234 15620 3240 15632
rect 2832 15592 3240 15620
rect 2832 15580 2838 15592
rect 3234 15580 3240 15592
rect 3292 15580 3298 15632
rect 7282 15620 7288 15632
rect 5368 15592 7288 15620
rect 3878 15512 3884 15564
rect 3936 15512 3942 15564
rect 4062 15512 4068 15564
rect 4120 15552 4126 15564
rect 4120 15524 4660 15552
rect 4120 15512 4126 15524
rect 198 15444 204 15496
rect 256 15484 262 15496
rect 3896 15484 3924 15512
rect 3973 15487 4031 15493
rect 3973 15484 3985 15487
rect 256 15456 3740 15484
rect 3896 15456 3985 15484
rect 256 15444 262 15456
rect 1394 15376 1400 15428
rect 1452 15416 1458 15428
rect 3602 15416 3608 15428
rect 1452 15388 3608 15416
rect 1452 15376 1458 15388
rect 3602 15376 3608 15388
rect 3660 15376 3666 15428
rect 3712 15416 3740 15456
rect 3973 15453 3985 15456
rect 4019 15453 4031 15487
rect 3973 15447 4031 15453
rect 4154 15444 4160 15496
rect 4212 15444 4218 15496
rect 4249 15487 4307 15493
rect 4249 15453 4261 15487
rect 4295 15484 4307 15487
rect 4338 15484 4344 15496
rect 4295 15456 4344 15484
rect 4295 15453 4307 15456
rect 4249 15447 4307 15453
rect 4338 15444 4344 15456
rect 4396 15444 4402 15496
rect 4632 15493 4660 15524
rect 4706 15512 4712 15564
rect 4764 15512 4770 15564
rect 4617 15487 4675 15493
rect 4617 15453 4629 15487
rect 4663 15484 4675 15487
rect 4890 15484 4896 15496
rect 4663 15456 4896 15484
rect 4663 15453 4675 15456
rect 4617 15447 4675 15453
rect 4890 15444 4896 15456
rect 4948 15444 4954 15496
rect 5166 15444 5172 15496
rect 5224 15444 5230 15496
rect 5261 15487 5319 15493
rect 5261 15453 5273 15487
rect 5307 15484 5319 15487
rect 5368 15484 5396 15592
rect 7282 15580 7288 15592
rect 7340 15580 7346 15632
rect 8312 15620 8340 15660
rect 8478 15648 8484 15700
rect 8536 15688 8542 15700
rect 8573 15691 8631 15697
rect 8573 15688 8585 15691
rect 8536 15660 8585 15688
rect 8536 15648 8542 15660
rect 8573 15657 8585 15660
rect 8619 15657 8631 15691
rect 9306 15688 9312 15700
rect 8573 15651 8631 15657
rect 8680 15660 9312 15688
rect 8680 15620 8708 15660
rect 9306 15648 9312 15660
rect 9364 15648 9370 15700
rect 9490 15648 9496 15700
rect 9548 15648 9554 15700
rect 10594 15648 10600 15700
rect 10652 15648 10658 15700
rect 10686 15648 10692 15700
rect 10744 15688 10750 15700
rect 16390 15688 16396 15700
rect 10744 15660 16396 15688
rect 10744 15648 10750 15660
rect 16390 15648 16396 15660
rect 16448 15648 16454 15700
rect 8312 15592 8708 15620
rect 8757 15623 8815 15629
rect 8757 15589 8769 15623
rect 8803 15620 8815 15623
rect 11146 15620 11152 15632
rect 8803 15592 11152 15620
rect 8803 15589 8815 15592
rect 8757 15583 8815 15589
rect 11146 15580 11152 15592
rect 11204 15580 11210 15632
rect 11808 15592 14780 15620
rect 6454 15512 6460 15564
rect 6512 15552 6518 15564
rect 7469 15555 7527 15561
rect 7469 15552 7481 15555
rect 6512 15524 7481 15552
rect 6512 15512 6518 15524
rect 7469 15521 7481 15524
rect 7515 15552 7527 15555
rect 11514 15552 11520 15564
rect 7515 15524 11520 15552
rect 7515 15521 7527 15524
rect 7469 15515 7527 15521
rect 11514 15512 11520 15524
rect 11572 15512 11578 15564
rect 6914 15484 6920 15496
rect 5307 15456 5396 15484
rect 5460 15456 6920 15484
rect 5307 15453 5319 15456
rect 5261 15447 5319 15453
rect 5460 15416 5488 15456
rect 6914 15444 6920 15456
rect 6972 15444 6978 15496
rect 7742 15484 7748 15496
rect 7392 15456 7748 15484
rect 3712 15388 3924 15416
rect 2406 15308 2412 15360
rect 2464 15348 2470 15360
rect 3789 15351 3847 15357
rect 3789 15348 3801 15351
rect 2464 15320 3801 15348
rect 2464 15308 2470 15320
rect 3789 15317 3801 15320
rect 3835 15317 3847 15351
rect 3896 15348 3924 15388
rect 4126 15388 5488 15416
rect 4126 15348 4154 15388
rect 6546 15376 6552 15428
rect 6604 15376 6610 15428
rect 3896 15320 4154 15348
rect 4985 15351 5043 15357
rect 3789 15311 3847 15317
rect 4985 15317 4997 15351
rect 5031 15348 5043 15351
rect 5442 15348 5448 15360
rect 5031 15320 5448 15348
rect 5031 15317 5043 15320
rect 4985 15311 5043 15317
rect 5442 15308 5448 15320
rect 5500 15308 5506 15360
rect 5534 15308 5540 15360
rect 5592 15348 5598 15360
rect 7392 15348 7420 15456
rect 7742 15444 7748 15456
rect 7800 15444 7806 15496
rect 8018 15444 8024 15496
rect 8076 15444 8082 15496
rect 8294 15444 8300 15496
rect 8352 15444 8358 15496
rect 8846 15444 8852 15496
rect 8904 15484 8910 15496
rect 8941 15487 8999 15493
rect 8941 15484 8953 15487
rect 8904 15456 8953 15484
rect 8904 15444 8910 15456
rect 8941 15453 8953 15456
rect 8987 15453 8999 15487
rect 8941 15447 8999 15453
rect 9030 15444 9036 15496
rect 9088 15444 9094 15496
rect 9217 15487 9275 15493
rect 9217 15453 9229 15487
rect 9263 15453 9275 15487
rect 9217 15447 9275 15453
rect 7834 15376 7840 15428
rect 7892 15416 7898 15428
rect 7929 15419 7987 15425
rect 7929 15416 7941 15419
rect 7892 15388 7941 15416
rect 7892 15376 7898 15388
rect 7929 15385 7941 15388
rect 7975 15385 7987 15419
rect 7929 15379 7987 15385
rect 8386 15376 8392 15428
rect 8444 15376 8450 15428
rect 9232 15416 9260 15447
rect 9306 15444 9312 15496
rect 9364 15444 9370 15496
rect 9508 15456 10364 15484
rect 9398 15416 9404 15428
rect 8496 15388 8708 15416
rect 9232 15388 9404 15416
rect 5592 15320 7420 15348
rect 5592 15308 5598 15320
rect 7466 15308 7472 15360
rect 7524 15348 7530 15360
rect 8496 15348 8524 15388
rect 7524 15320 8524 15348
rect 7524 15308 7530 15320
rect 8570 15308 8576 15360
rect 8628 15357 8634 15360
rect 8628 15351 8647 15357
rect 8635 15317 8647 15351
rect 8680 15348 8708 15388
rect 9398 15376 9404 15388
rect 9456 15376 9462 15428
rect 9508 15348 9536 15456
rect 10336 15416 10364 15456
rect 10410 15444 10416 15496
rect 10468 15484 10474 15496
rect 10594 15484 10600 15496
rect 10468 15456 10600 15484
rect 10468 15444 10474 15456
rect 10594 15444 10600 15456
rect 10652 15444 10658 15496
rect 11054 15444 11060 15496
rect 11112 15444 11118 15496
rect 11422 15444 11428 15496
rect 11480 15444 11486 15496
rect 11698 15444 11704 15496
rect 11756 15444 11762 15496
rect 11808 15416 11836 15592
rect 12618 15512 12624 15564
rect 12676 15512 12682 15564
rect 12710 15512 12716 15564
rect 12768 15552 12774 15564
rect 14752 15552 14780 15592
rect 14826 15580 14832 15632
rect 14884 15580 14890 15632
rect 16758 15552 16764 15564
rect 12768 15524 13400 15552
rect 14752 15524 16764 15552
rect 12768 15512 12774 15524
rect 12529 15487 12587 15493
rect 12529 15453 12541 15487
rect 12575 15484 12587 15487
rect 12575 15456 12756 15484
rect 12575 15453 12587 15456
rect 12529 15447 12587 15453
rect 10336 15388 11836 15416
rect 12342 15376 12348 15428
rect 12400 15416 12406 15428
rect 12437 15419 12495 15425
rect 12437 15416 12449 15419
rect 12400 15388 12449 15416
rect 12400 15376 12406 15388
rect 12437 15385 12449 15388
rect 12483 15416 12495 15419
rect 12618 15416 12624 15428
rect 12483 15388 12624 15416
rect 12483 15385 12495 15388
rect 12437 15379 12495 15385
rect 12618 15376 12624 15388
rect 12676 15376 12682 15428
rect 12728 15416 12756 15456
rect 12802 15444 12808 15496
rect 12860 15444 12866 15496
rect 13372 15493 13400 15524
rect 16758 15512 16764 15524
rect 16816 15512 16822 15564
rect 13357 15487 13415 15493
rect 13357 15453 13369 15487
rect 13403 15453 13415 15487
rect 13357 15447 13415 15453
rect 12986 15416 12992 15428
rect 12728 15388 12992 15416
rect 12986 15376 12992 15388
rect 13044 15376 13050 15428
rect 13372 15416 13400 15447
rect 15010 15444 15016 15496
rect 15068 15444 15074 15496
rect 15289 15487 15347 15493
rect 15289 15453 15301 15487
rect 15335 15453 15347 15487
rect 15289 15447 15347 15453
rect 15304 15416 15332 15447
rect 13372 15388 15332 15416
rect 8680 15320 9536 15348
rect 8628 15311 8647 15317
rect 8628 15308 8634 15311
rect 9766 15308 9772 15360
rect 9824 15348 9830 15360
rect 10962 15348 10968 15360
rect 9824 15320 10968 15348
rect 9824 15308 9830 15320
rect 10962 15308 10968 15320
rect 11020 15308 11026 15360
rect 11514 15308 11520 15360
rect 11572 15348 11578 15360
rect 13173 15351 13231 15357
rect 13173 15348 13185 15351
rect 11572 15320 13185 15348
rect 11572 15308 11578 15320
rect 13173 15317 13185 15320
rect 13219 15317 13231 15351
rect 13173 15311 13231 15317
rect 15194 15308 15200 15360
rect 15252 15308 15258 15360
rect 1104 15258 18860 15280
rect 1104 15206 2610 15258
rect 2662 15206 2674 15258
rect 2726 15206 2738 15258
rect 2790 15206 2802 15258
rect 2854 15206 2866 15258
rect 2918 15206 7610 15258
rect 7662 15206 7674 15258
rect 7726 15206 7738 15258
rect 7790 15206 7802 15258
rect 7854 15206 7866 15258
rect 7918 15206 12610 15258
rect 12662 15206 12674 15258
rect 12726 15206 12738 15258
rect 12790 15206 12802 15258
rect 12854 15206 12866 15258
rect 12918 15206 17610 15258
rect 17662 15206 17674 15258
rect 17726 15206 17738 15258
rect 17790 15206 17802 15258
rect 17854 15206 17866 15258
rect 17918 15206 18860 15258
rect 1104 15184 18860 15206
rect 1302 15104 1308 15156
rect 1360 15144 1366 15156
rect 1765 15147 1823 15153
rect 1765 15144 1777 15147
rect 1360 15116 1777 15144
rect 1360 15104 1366 15116
rect 1765 15113 1777 15116
rect 1811 15113 1823 15147
rect 1765 15107 1823 15113
rect 8202 15104 8208 15156
rect 8260 15144 8266 15156
rect 9766 15144 9772 15156
rect 8260 15116 9772 15144
rect 8260 15104 8266 15116
rect 9766 15104 9772 15116
rect 9824 15104 9830 15156
rect 9950 15104 9956 15156
rect 10008 15144 10014 15156
rect 10008 15116 14145 15144
rect 10008 15104 10014 15116
rect 1118 15036 1124 15088
rect 1176 15076 1182 15088
rect 1176 15048 1900 15076
rect 1176 15036 1182 15048
rect 1872 15017 1900 15048
rect 5258 15036 5264 15088
rect 5316 15036 5322 15088
rect 8018 15036 8024 15088
rect 8076 15076 8082 15088
rect 8076 15048 10916 15076
rect 8076 15036 8082 15048
rect 1581 15011 1639 15017
rect 1581 14977 1593 15011
rect 1627 14977 1639 15011
rect 1581 14971 1639 14977
rect 1857 15011 1915 15017
rect 1857 14977 1869 15011
rect 1903 14977 1915 15011
rect 1857 14971 1915 14977
rect 1596 14940 1624 14971
rect 4522 14968 4528 15020
rect 4580 14968 4586 15020
rect 4614 14968 4620 15020
rect 4672 14968 4678 15020
rect 4801 15011 4859 15017
rect 4801 14977 4813 15011
rect 4847 15008 4859 15011
rect 8386 15008 8392 15020
rect 4847 14980 8392 15008
rect 4847 14977 4859 14980
rect 4801 14971 4859 14977
rect 1762 14940 1768 14952
rect 1596 14912 1768 14940
rect 1762 14900 1768 14912
rect 1820 14940 1826 14952
rect 2314 14940 2320 14952
rect 1820 14912 2320 14940
rect 1820 14900 1826 14912
rect 2314 14900 2320 14912
rect 2372 14900 2378 14952
rect 3878 14900 3884 14952
rect 3936 14940 3942 14952
rect 4816 14940 4844 14971
rect 8386 14968 8392 14980
rect 8444 14968 8450 15020
rect 9585 15011 9643 15017
rect 9585 14977 9597 15011
rect 9631 15008 9643 15011
rect 9766 15008 9772 15020
rect 9631 14980 9772 15008
rect 9631 14977 9643 14980
rect 9585 14971 9643 14977
rect 9766 14968 9772 14980
rect 9824 14968 9830 15020
rect 10134 14968 10140 15020
rect 10192 14968 10198 15020
rect 10226 14968 10232 15020
rect 10284 15008 10290 15020
rect 10781 15011 10839 15017
rect 10781 15008 10793 15011
rect 10284 14980 10793 15008
rect 10284 14968 10290 14980
rect 10781 14977 10793 14980
rect 10827 14977 10839 15011
rect 10781 14971 10839 14977
rect 8478 14940 8484 14952
rect 3936 14912 4844 14940
rect 5506 14912 8484 14940
rect 3936 14900 3942 14912
rect 1397 14875 1455 14881
rect 1397 14841 1409 14875
rect 1443 14872 1455 14875
rect 3970 14872 3976 14884
rect 1443 14844 3976 14872
rect 1443 14841 1455 14844
rect 1397 14835 1455 14841
rect 3970 14832 3976 14844
rect 4028 14832 4034 14884
rect 5506 14872 5534 14912
rect 8478 14900 8484 14912
rect 8536 14900 8542 14952
rect 8570 14900 8576 14952
rect 8628 14940 8634 14952
rect 9306 14940 9312 14952
rect 8628 14912 9312 14940
rect 8628 14900 8634 14912
rect 9306 14900 9312 14912
rect 9364 14900 9370 14952
rect 9674 14900 9680 14952
rect 9732 14900 9738 14952
rect 10321 14943 10379 14949
rect 10321 14909 10333 14943
rect 10367 14940 10379 14943
rect 10410 14940 10416 14952
rect 10367 14912 10416 14940
rect 10367 14909 10379 14912
rect 10321 14903 10379 14909
rect 10410 14900 10416 14912
rect 10468 14900 10474 14952
rect 10689 14943 10747 14949
rect 10689 14909 10701 14943
rect 10735 14909 10747 14943
rect 10888 14940 10916 15048
rect 11238 15036 11244 15088
rect 11296 15076 11302 15088
rect 11885 15079 11943 15085
rect 11885 15076 11897 15079
rect 11296 15048 11897 15076
rect 11296 15036 11302 15048
rect 11885 15045 11897 15048
rect 11931 15045 11943 15079
rect 12802 15076 12808 15088
rect 11885 15039 11943 15045
rect 12176 15048 12808 15076
rect 11701 15011 11759 15017
rect 11701 14977 11713 15011
rect 11747 15008 11759 15011
rect 12176 15008 12204 15048
rect 12802 15036 12808 15048
rect 12860 15036 12866 15088
rect 13722 15076 13728 15088
rect 13004 15048 13728 15076
rect 11747 14980 12204 15008
rect 12345 15011 12403 15017
rect 11747 14977 11759 14980
rect 11701 14971 11759 14977
rect 12345 14977 12357 15011
rect 12391 14977 12403 15011
rect 12345 14971 12403 14977
rect 12360 14940 12388 14971
rect 12434 14968 12440 15020
rect 12492 15008 12498 15020
rect 12529 15011 12587 15017
rect 12529 15008 12541 15011
rect 12492 14980 12541 15008
rect 12492 14968 12498 14980
rect 12529 14977 12541 14980
rect 12575 14977 12587 15011
rect 12529 14971 12587 14977
rect 12894 14968 12900 15020
rect 12952 14968 12958 15020
rect 13004 15017 13032 15048
rect 13722 15036 13728 15048
rect 13780 15036 13786 15088
rect 12989 15011 13047 15017
rect 12989 14977 13001 15011
rect 13035 14977 13047 15011
rect 12989 14971 13047 14977
rect 13265 15011 13323 15017
rect 13265 14977 13277 15011
rect 13311 14977 13323 15011
rect 13265 14971 13323 14977
rect 13078 14940 13084 14952
rect 10888 14912 13084 14940
rect 10689 14903 10747 14909
rect 4080 14844 5534 14872
rect 3234 14764 3240 14816
rect 3292 14804 3298 14816
rect 4080 14804 4108 14844
rect 5626 14832 5632 14884
rect 5684 14872 5690 14884
rect 10704 14872 10732 14903
rect 13078 14900 13084 14912
rect 13136 14900 13142 14952
rect 13280 14940 13308 14971
rect 13354 14968 13360 15020
rect 13412 14968 13418 15020
rect 13446 14968 13452 15020
rect 13504 15008 13510 15020
rect 13541 15011 13599 15017
rect 13541 15008 13553 15011
rect 13504 14980 13553 15008
rect 13504 14968 13510 14980
rect 13541 14977 13553 14980
rect 13587 14977 13599 15011
rect 13541 14971 13599 14977
rect 13814 14968 13820 15020
rect 13872 15008 13878 15020
rect 14117 15017 14145 15116
rect 14274 15036 14280 15088
rect 14332 15076 14338 15088
rect 14332 15048 17632 15076
rect 14332 15036 14338 15048
rect 13909 15011 13967 15017
rect 13909 15008 13921 15011
rect 13872 14980 13921 15008
rect 13872 14968 13878 14980
rect 13909 14977 13921 14980
rect 13955 14977 13967 15011
rect 13909 14971 13967 14977
rect 14102 15011 14160 15017
rect 14102 14977 14114 15011
rect 14148 14977 14160 15011
rect 14102 14971 14160 14977
rect 16666 14968 16672 15020
rect 16724 14968 16730 15020
rect 17129 15011 17187 15017
rect 17129 14977 17141 15011
rect 17175 14977 17187 15011
rect 17129 14971 17187 14977
rect 13280 14912 14688 14940
rect 5684 14844 10732 14872
rect 5684 14832 5690 14844
rect 11146 14832 11152 14884
rect 11204 14872 11210 14884
rect 12618 14872 12624 14884
rect 11204 14844 12624 14872
rect 11204 14832 11210 14844
rect 12618 14832 12624 14844
rect 12676 14832 12682 14884
rect 12897 14875 12955 14881
rect 12897 14841 12909 14875
rect 12943 14872 12955 14875
rect 13170 14872 13176 14884
rect 12943 14844 13176 14872
rect 12943 14841 12955 14844
rect 12897 14835 12955 14841
rect 13170 14832 13176 14844
rect 13228 14832 13234 14884
rect 14660 14872 14688 14912
rect 14734 14900 14740 14952
rect 14792 14900 14798 14952
rect 16022 14900 16028 14952
rect 16080 14940 16086 14952
rect 17144 14940 17172 14971
rect 17402 14968 17408 15020
rect 17460 14968 17466 15020
rect 17604 14949 17632 15048
rect 18138 14968 18144 15020
rect 18196 14968 18202 15020
rect 16080 14912 17172 14940
rect 17589 14943 17647 14949
rect 16080 14900 16086 14912
rect 17589 14909 17601 14943
rect 17635 14909 17647 14943
rect 17589 14903 17647 14909
rect 15102 14872 15108 14884
rect 14660 14844 15108 14872
rect 15102 14832 15108 14844
rect 15160 14832 15166 14884
rect 3292 14776 4108 14804
rect 3292 14764 3298 14776
rect 8478 14764 8484 14816
rect 8536 14804 8542 14816
rect 9490 14804 9496 14816
rect 8536 14776 9496 14804
rect 8536 14764 8542 14776
rect 9490 14764 9496 14776
rect 9548 14764 9554 14816
rect 10594 14764 10600 14816
rect 10652 14804 10658 14816
rect 10965 14807 11023 14813
rect 10965 14804 10977 14807
rect 10652 14776 10977 14804
rect 10652 14764 10658 14776
rect 10965 14773 10977 14776
rect 11011 14773 11023 14807
rect 10965 14767 11023 14773
rect 11514 14764 11520 14816
rect 11572 14764 11578 14816
rect 11698 14764 11704 14816
rect 11756 14804 11762 14816
rect 15194 14804 15200 14816
rect 11756 14776 15200 14804
rect 11756 14764 11762 14776
rect 15194 14764 15200 14776
rect 15252 14764 15258 14816
rect 1104 14714 18860 14736
rect 1104 14662 1950 14714
rect 2002 14662 2014 14714
rect 2066 14662 2078 14714
rect 2130 14662 2142 14714
rect 2194 14662 2206 14714
rect 2258 14662 6950 14714
rect 7002 14662 7014 14714
rect 7066 14662 7078 14714
rect 7130 14662 7142 14714
rect 7194 14662 7206 14714
rect 7258 14662 11950 14714
rect 12002 14662 12014 14714
rect 12066 14662 12078 14714
rect 12130 14662 12142 14714
rect 12194 14662 12206 14714
rect 12258 14662 16950 14714
rect 17002 14662 17014 14714
rect 17066 14662 17078 14714
rect 17130 14662 17142 14714
rect 17194 14662 17206 14714
rect 17258 14662 18860 14714
rect 1104 14640 18860 14662
rect 1762 14560 1768 14612
rect 1820 14560 1826 14612
rect 2222 14560 2228 14612
rect 2280 14600 2286 14612
rect 6178 14600 6184 14612
rect 2280 14572 6184 14600
rect 2280 14560 2286 14572
rect 6178 14560 6184 14572
rect 6236 14560 6242 14612
rect 8386 14560 8392 14612
rect 8444 14600 8450 14612
rect 8444 14572 9444 14600
rect 8444 14560 8450 14572
rect 6546 14492 6552 14544
rect 6604 14532 6610 14544
rect 8570 14532 8576 14544
rect 6604 14504 8576 14532
rect 6604 14492 6610 14504
rect 8570 14492 8576 14504
rect 8628 14492 8634 14544
rect 8754 14492 8760 14544
rect 8812 14532 8818 14544
rect 9416 14532 9444 14572
rect 9490 14560 9496 14612
rect 9548 14600 9554 14612
rect 9585 14603 9643 14609
rect 9585 14600 9597 14603
rect 9548 14572 9597 14600
rect 9548 14560 9554 14572
rect 9585 14569 9597 14572
rect 9631 14600 9643 14603
rect 10686 14600 10692 14612
rect 9631 14572 10692 14600
rect 9631 14569 9643 14572
rect 9585 14563 9643 14569
rect 10686 14560 10692 14572
rect 10744 14560 10750 14612
rect 10962 14560 10968 14612
rect 11020 14600 11026 14612
rect 11882 14600 11888 14612
rect 11020 14572 11888 14600
rect 11020 14560 11026 14572
rect 11882 14560 11888 14572
rect 11940 14560 11946 14612
rect 12250 14560 12256 14612
rect 12308 14600 12314 14612
rect 12618 14600 12624 14612
rect 12308 14572 12624 14600
rect 12308 14560 12314 14572
rect 12618 14560 12624 14572
rect 12676 14560 12682 14612
rect 12710 14560 12716 14612
rect 12768 14600 12774 14612
rect 14090 14600 14096 14612
rect 12768 14572 14096 14600
rect 12768 14560 12774 14572
rect 14090 14560 14096 14572
rect 14148 14560 14154 14612
rect 15746 14560 15752 14612
rect 15804 14600 15810 14612
rect 16393 14603 16451 14609
rect 16393 14600 16405 14603
rect 15804 14572 16405 14600
rect 15804 14560 15810 14572
rect 16393 14569 16405 14572
rect 16439 14569 16451 14603
rect 16393 14563 16451 14569
rect 16482 14560 16488 14612
rect 16540 14600 16546 14612
rect 16540 14572 17724 14600
rect 16540 14560 16546 14572
rect 11146 14532 11152 14544
rect 8812 14504 9352 14532
rect 9416 14504 11152 14532
rect 8812 14492 8818 14504
rect 9324 14476 9352 14504
rect 11146 14492 11152 14504
rect 11204 14492 11210 14544
rect 11238 14492 11244 14544
rect 11296 14532 11302 14544
rect 11698 14532 11704 14544
rect 11296 14504 11704 14532
rect 11296 14492 11302 14504
rect 11698 14492 11704 14504
rect 11756 14492 11762 14544
rect 11808 14504 12848 14532
rect 1670 14424 1676 14476
rect 1728 14464 1734 14476
rect 1854 14464 1860 14476
rect 1728 14436 1860 14464
rect 1728 14424 1734 14436
rect 1854 14424 1860 14436
rect 1912 14464 1918 14476
rect 2041 14467 2099 14473
rect 2041 14464 2053 14467
rect 1912 14436 2053 14464
rect 1912 14424 1918 14436
rect 2041 14433 2053 14436
rect 2087 14433 2099 14467
rect 2041 14427 2099 14433
rect 2222 14424 2228 14476
rect 2280 14424 2286 14476
rect 2958 14424 2964 14476
rect 3016 14464 3022 14476
rect 5994 14464 6000 14476
rect 3016 14436 6000 14464
rect 3016 14424 3022 14436
rect 5994 14424 6000 14436
rect 6052 14424 6058 14476
rect 6472 14436 8064 14464
rect 1946 14356 1952 14408
rect 2004 14356 2010 14408
rect 2130 14356 2136 14408
rect 2188 14356 2194 14408
rect 4706 14356 4712 14408
rect 4764 14356 4770 14408
rect 4982 14356 4988 14408
rect 5040 14396 5046 14408
rect 5166 14396 5172 14408
rect 5040 14368 5172 14396
rect 5040 14356 5046 14368
rect 5166 14356 5172 14368
rect 5224 14356 5230 14408
rect 5258 14356 5264 14408
rect 5316 14396 5322 14408
rect 6472 14396 6500 14436
rect 5316 14368 6500 14396
rect 8036 14396 8064 14436
rect 9122 14424 9128 14476
rect 9180 14464 9186 14476
rect 9217 14467 9275 14473
rect 9217 14464 9229 14467
rect 9180 14436 9229 14464
rect 9180 14424 9186 14436
rect 9217 14433 9229 14436
rect 9263 14433 9275 14467
rect 9217 14427 9275 14433
rect 9306 14424 9312 14476
rect 9364 14464 9370 14476
rect 11808 14464 11836 14504
rect 9364 14436 11836 14464
rect 12820 14464 12848 14504
rect 12986 14492 12992 14544
rect 13044 14532 13050 14544
rect 13354 14532 13360 14544
rect 13044 14504 13360 14532
rect 13044 14492 13050 14504
rect 13354 14492 13360 14504
rect 13412 14492 13418 14544
rect 13630 14492 13636 14544
rect 13688 14532 13694 14544
rect 16945 14535 17003 14541
rect 13688 14504 16804 14532
rect 13688 14492 13694 14504
rect 12820 14436 13400 14464
rect 9364 14424 9370 14436
rect 12716 14408 12768 14414
rect 8036 14368 10640 14396
rect 5316 14356 5322 14368
rect 3602 14288 3608 14340
rect 3660 14328 3666 14340
rect 9585 14331 9643 14337
rect 9585 14328 9597 14331
rect 3660 14300 9597 14328
rect 3660 14288 3666 14300
rect 9585 14297 9597 14300
rect 9631 14297 9643 14331
rect 10502 14328 10508 14340
rect 9585 14291 9643 14297
rect 9692 14300 10508 14328
rect 4890 14220 4896 14272
rect 4948 14220 4954 14272
rect 5902 14220 5908 14272
rect 5960 14260 5966 14272
rect 9692 14260 9720 14300
rect 10502 14288 10508 14300
rect 10560 14288 10566 14340
rect 10612 14328 10640 14368
rect 10686 14356 10692 14408
rect 10744 14396 10750 14408
rect 11701 14399 11759 14405
rect 11701 14396 11713 14399
rect 10744 14368 11713 14396
rect 10744 14356 10750 14368
rect 11701 14365 11713 14368
rect 11747 14365 11759 14399
rect 12069 14399 12127 14405
rect 12069 14396 12081 14399
rect 11701 14359 11759 14365
rect 11808 14368 12081 14396
rect 11808 14328 11836 14368
rect 12069 14365 12081 14368
rect 12115 14365 12127 14399
rect 12069 14359 12127 14365
rect 12986 14356 12992 14408
rect 13044 14396 13050 14408
rect 13372 14405 13400 14436
rect 13446 14424 13452 14476
rect 13504 14464 13510 14476
rect 13504 14436 14596 14464
rect 13504 14424 13510 14436
rect 13173 14399 13231 14405
rect 13044 14368 13124 14396
rect 13044 14356 13050 14368
rect 12716 14350 12768 14356
rect 10612 14300 11836 14328
rect 11882 14288 11888 14340
rect 11940 14288 11946 14340
rect 13096 14337 13124 14368
rect 13173 14365 13185 14399
rect 13219 14365 13231 14399
rect 13173 14359 13231 14365
rect 13357 14399 13415 14405
rect 13357 14365 13369 14399
rect 13403 14365 13415 14399
rect 13357 14359 13415 14365
rect 13081 14331 13139 14337
rect 13081 14297 13093 14331
rect 13127 14297 13139 14331
rect 13188 14328 13216 14359
rect 13906 14356 13912 14408
rect 13964 14396 13970 14408
rect 14093 14399 14151 14405
rect 14093 14396 14105 14399
rect 13964 14368 14105 14396
rect 13964 14356 13970 14368
rect 14093 14365 14105 14368
rect 14139 14365 14151 14399
rect 14093 14359 14151 14365
rect 14274 14356 14280 14408
rect 14332 14356 14338 14408
rect 14568 14405 14596 14436
rect 15930 14424 15936 14476
rect 15988 14464 15994 14476
rect 16482 14464 16488 14476
rect 15988 14436 16488 14464
rect 15988 14424 15994 14436
rect 16482 14424 16488 14436
rect 16540 14424 16546 14476
rect 14553 14399 14611 14405
rect 14553 14365 14565 14399
rect 14599 14365 14611 14399
rect 14553 14359 14611 14365
rect 16117 14399 16175 14405
rect 16117 14365 16129 14399
rect 16163 14396 16175 14399
rect 16390 14396 16396 14408
rect 16163 14368 16396 14396
rect 16163 14365 16175 14368
rect 16117 14359 16175 14365
rect 16390 14356 16396 14368
rect 16448 14356 16454 14408
rect 16666 14356 16672 14408
rect 16724 14356 16730 14408
rect 16776 14405 16804 14504
rect 16945 14501 16957 14535
rect 16991 14532 17003 14535
rect 17494 14532 17500 14544
rect 16991 14504 17500 14532
rect 16991 14501 17003 14504
rect 16945 14495 17003 14501
rect 17494 14492 17500 14504
rect 17552 14492 17558 14544
rect 17696 14541 17724 14572
rect 17681 14535 17739 14541
rect 17681 14501 17693 14535
rect 17727 14501 17739 14535
rect 17681 14495 17739 14501
rect 16761 14399 16819 14405
rect 16761 14365 16773 14399
rect 16807 14365 16819 14399
rect 18230 14396 18236 14408
rect 16761 14359 16819 14365
rect 16868 14368 18236 14396
rect 13538 14328 13544 14340
rect 13188 14300 13544 14328
rect 13081 14291 13139 14297
rect 13538 14288 13544 14300
rect 13596 14288 13602 14340
rect 14182 14288 14188 14340
rect 14240 14288 14246 14340
rect 16577 14331 16635 14337
rect 15304 14300 16528 14328
rect 5960 14232 9720 14260
rect 5960 14220 5966 14232
rect 9766 14220 9772 14272
rect 9824 14220 9830 14272
rect 10962 14220 10968 14272
rect 11020 14260 11026 14272
rect 11333 14263 11391 14269
rect 11333 14260 11345 14263
rect 11020 14232 11345 14260
rect 11020 14220 11026 14232
rect 11333 14229 11345 14232
rect 11379 14229 11391 14263
rect 11333 14223 11391 14229
rect 11514 14220 11520 14272
rect 11572 14220 11578 14272
rect 11609 14263 11667 14269
rect 11609 14229 11621 14263
rect 11655 14260 11667 14263
rect 11974 14260 11980 14272
rect 11655 14232 11980 14260
rect 11655 14229 11667 14232
rect 11609 14223 11667 14229
rect 11974 14220 11980 14232
rect 12032 14260 12038 14272
rect 12434 14260 12440 14272
rect 12032 14232 12440 14260
rect 12032 14220 12038 14232
rect 12434 14220 12440 14232
rect 12492 14220 12498 14272
rect 13357 14263 13415 14269
rect 13357 14229 13369 14263
rect 13403 14260 13415 14263
rect 15304 14260 15332 14300
rect 13403 14232 15332 14260
rect 13403 14229 13415 14232
rect 13357 14223 13415 14229
rect 16298 14220 16304 14272
rect 16356 14260 16362 14272
rect 16393 14263 16451 14269
rect 16393 14260 16405 14263
rect 16356 14232 16405 14260
rect 16356 14220 16362 14232
rect 16393 14229 16405 14232
rect 16439 14229 16451 14263
rect 16500 14260 16528 14300
rect 16577 14297 16589 14331
rect 16623 14328 16635 14331
rect 16868 14328 16896 14368
rect 18230 14356 18236 14368
rect 18288 14356 18294 14408
rect 16623 14300 16896 14328
rect 16945 14331 17003 14337
rect 16623 14297 16635 14300
rect 16577 14291 16635 14297
rect 16945 14297 16957 14331
rect 16991 14328 17003 14331
rect 16991 14300 18000 14328
rect 16991 14297 17003 14300
rect 16945 14291 17003 14297
rect 16666 14260 16672 14272
rect 16500 14232 16672 14260
rect 16393 14223 16451 14229
rect 16666 14220 16672 14232
rect 16724 14220 16730 14272
rect 16758 14220 16764 14272
rect 16816 14260 16822 14272
rect 16960 14260 16988 14291
rect 16816 14232 16988 14260
rect 16816 14220 16822 14232
rect 17126 14220 17132 14272
rect 17184 14260 17190 14272
rect 17589 14263 17647 14269
rect 17589 14260 17601 14263
rect 17184 14232 17601 14260
rect 17184 14220 17190 14232
rect 17589 14229 17601 14232
rect 17635 14229 17647 14263
rect 17972 14260 18000 14300
rect 18046 14288 18052 14340
rect 18104 14288 18110 14340
rect 18874 14260 18880 14272
rect 17972 14232 18880 14260
rect 17589 14223 17647 14229
rect 18874 14220 18880 14232
rect 18932 14220 18938 14272
rect 1104 14170 18860 14192
rect 1104 14118 2610 14170
rect 2662 14118 2674 14170
rect 2726 14118 2738 14170
rect 2790 14118 2802 14170
rect 2854 14118 2866 14170
rect 2918 14118 7610 14170
rect 7662 14118 7674 14170
rect 7726 14118 7738 14170
rect 7790 14118 7802 14170
rect 7854 14118 7866 14170
rect 7918 14118 12610 14170
rect 12662 14118 12674 14170
rect 12726 14118 12738 14170
rect 12790 14118 12802 14170
rect 12854 14118 12866 14170
rect 12918 14118 17610 14170
rect 17662 14118 17674 14170
rect 17726 14118 17738 14170
rect 17790 14118 17802 14170
rect 17854 14118 17866 14170
rect 17918 14118 18860 14170
rect 1104 14096 18860 14118
rect 2866 14016 2872 14068
rect 2924 14056 2930 14068
rect 3234 14056 3240 14068
rect 2924 14028 3240 14056
rect 2924 14016 2930 14028
rect 3234 14016 3240 14028
rect 3292 14016 3298 14068
rect 4614 14016 4620 14068
rect 4672 14056 4678 14068
rect 7469 14059 7527 14065
rect 7469 14056 7481 14059
rect 4672 14028 7481 14056
rect 4672 14016 4678 14028
rect 7469 14025 7481 14028
rect 7515 14025 7527 14059
rect 7469 14019 7527 14025
rect 8573 14059 8631 14065
rect 8573 14025 8585 14059
rect 8619 14056 8631 14059
rect 8662 14056 8668 14068
rect 8619 14028 8668 14056
rect 8619 14025 8631 14028
rect 8573 14019 8631 14025
rect 8662 14016 8668 14028
rect 8720 14016 8726 14068
rect 9214 14016 9220 14068
rect 9272 14016 9278 14068
rect 9306 14016 9312 14068
rect 9364 14016 9370 14068
rect 11146 14016 11152 14068
rect 11204 14056 11210 14068
rect 13630 14056 13636 14068
rect 11204 14028 13636 14056
rect 11204 14016 11210 14028
rect 13630 14016 13636 14028
rect 13688 14016 13694 14068
rect 13814 14016 13820 14068
rect 13872 14056 13878 14068
rect 16022 14056 16028 14068
rect 13872 14028 16028 14056
rect 13872 14016 13878 14028
rect 16022 14016 16028 14028
rect 16080 14016 16086 14068
rect 3418 13988 3424 14000
rect 2746 13960 3424 13988
rect 1486 13880 1492 13932
rect 1544 13880 1550 13932
rect 2746 13929 2774 13960
rect 3418 13948 3424 13960
rect 3476 13948 3482 14000
rect 5261 13991 5319 13997
rect 5261 13957 5273 13991
rect 5307 13988 5319 13991
rect 5350 13988 5356 14000
rect 5307 13960 5356 13988
rect 5307 13957 5319 13960
rect 5261 13951 5319 13957
rect 5350 13948 5356 13960
rect 5408 13988 5414 14000
rect 7285 13991 7343 13997
rect 7285 13988 7297 13991
rect 5408 13960 5948 13988
rect 5408 13948 5414 13960
rect 5920 13932 5948 13960
rect 6012 13960 7297 13988
rect 2705 13923 2774 13929
rect 2705 13889 2717 13923
rect 2751 13892 2774 13923
rect 2751 13889 2763 13892
rect 2705 13883 2763 13889
rect 2866 13880 2872 13932
rect 2924 13880 2930 13932
rect 2958 13880 2964 13932
rect 3016 13880 3022 13932
rect 3053 13923 3111 13929
rect 3053 13889 3065 13923
rect 3099 13920 3111 13923
rect 3878 13920 3884 13932
rect 3099 13892 3884 13920
rect 3099 13889 3111 13892
rect 3053 13883 3111 13889
rect 3878 13880 3884 13892
rect 3936 13880 3942 13932
rect 4798 13880 4804 13932
rect 4856 13920 4862 13932
rect 5718 13920 5724 13932
rect 4856 13892 5724 13920
rect 4856 13880 4862 13892
rect 5718 13880 5724 13892
rect 5776 13880 5782 13932
rect 5902 13880 5908 13932
rect 5960 13880 5966 13932
rect 1765 13855 1823 13861
rect 1765 13821 1777 13855
rect 1811 13852 1823 13855
rect 3234 13852 3240 13864
rect 1811 13824 3240 13852
rect 1811 13821 1823 13824
rect 1765 13815 1823 13821
rect 3234 13812 3240 13824
rect 3292 13812 3298 13864
rect 5166 13852 5172 13864
rect 4816 13824 5172 13852
rect 290 13744 296 13796
rect 348 13784 354 13796
rect 4816 13784 4844 13824
rect 5166 13812 5172 13824
rect 5224 13812 5230 13864
rect 5350 13812 5356 13864
rect 5408 13852 5414 13864
rect 5534 13852 5540 13864
rect 5408 13824 5540 13852
rect 5408 13812 5414 13824
rect 5534 13812 5540 13824
rect 5592 13852 5598 13864
rect 5629 13855 5687 13861
rect 5629 13852 5641 13855
rect 5592 13824 5641 13852
rect 5592 13812 5598 13824
rect 5629 13821 5641 13824
rect 5675 13821 5687 13855
rect 5629 13815 5687 13821
rect 5810 13812 5816 13864
rect 5868 13852 5874 13864
rect 6012 13852 6040 13960
rect 7285 13957 7297 13960
rect 7331 13957 7343 13991
rect 7285 13951 7343 13957
rect 7653 13991 7711 13997
rect 7653 13957 7665 13991
rect 7699 13988 7711 13991
rect 8110 13988 8116 14000
rect 7699 13960 8116 13988
rect 7699 13957 7711 13960
rect 7653 13951 7711 13957
rect 8110 13948 8116 13960
rect 8168 13948 8174 14000
rect 9324 13988 9352 14016
rect 9324 13960 13032 13988
rect 6089 13923 6147 13929
rect 6089 13889 6101 13923
rect 6135 13920 6147 13923
rect 6362 13920 6368 13932
rect 6135 13892 6368 13920
rect 6135 13889 6147 13892
rect 6089 13883 6147 13889
rect 6362 13880 6368 13892
rect 6420 13880 6426 13932
rect 6454 13880 6460 13932
rect 6512 13880 6518 13932
rect 6638 13880 6644 13932
rect 6696 13880 6702 13932
rect 6825 13923 6883 13929
rect 6825 13889 6837 13923
rect 6871 13920 6883 13923
rect 7742 13920 7748 13932
rect 6871 13892 7748 13920
rect 6871 13889 6883 13892
rect 6825 13883 6883 13889
rect 7742 13880 7748 13892
rect 7800 13880 7806 13932
rect 7837 13923 7895 13929
rect 7837 13889 7849 13923
rect 7883 13920 7895 13923
rect 8018 13920 8024 13932
rect 7883 13892 8024 13920
rect 7883 13889 7895 13892
rect 7837 13883 7895 13889
rect 8018 13880 8024 13892
rect 8076 13880 8082 13932
rect 8662 13880 8668 13932
rect 8720 13920 8726 13932
rect 8757 13923 8815 13929
rect 8757 13920 8769 13923
rect 8720 13892 8769 13920
rect 8720 13880 8726 13892
rect 8757 13889 8769 13892
rect 8803 13889 8815 13923
rect 8757 13883 8815 13889
rect 8849 13923 8907 13929
rect 8849 13889 8861 13923
rect 8895 13889 8907 13923
rect 8849 13883 8907 13889
rect 5868 13824 6040 13852
rect 6181 13855 6239 13861
rect 5868 13812 5874 13824
rect 6181 13821 6193 13855
rect 6227 13852 6239 13855
rect 6472 13852 6500 13880
rect 8478 13852 8484 13864
rect 6227 13824 6500 13852
rect 6656 13824 8484 13852
rect 6227 13821 6239 13824
rect 6181 13815 6239 13821
rect 348 13756 4844 13784
rect 348 13744 354 13756
rect 4982 13744 4988 13796
rect 5040 13784 5046 13796
rect 6656 13784 6684 13824
rect 8478 13812 8484 13824
rect 8536 13852 8542 13864
rect 8573 13855 8631 13861
rect 8573 13852 8585 13855
rect 8536 13824 8585 13852
rect 8536 13812 8542 13824
rect 8573 13821 8585 13824
rect 8619 13821 8631 13855
rect 8864 13852 8892 13883
rect 8938 13880 8944 13932
rect 8996 13880 9002 13932
rect 9306 13880 9312 13932
rect 9364 13920 9370 13932
rect 12161 13923 12219 13929
rect 12161 13920 12173 13923
rect 9364 13892 12173 13920
rect 9364 13880 9370 13892
rect 12161 13889 12173 13892
rect 12207 13889 12219 13923
rect 12161 13883 12219 13889
rect 12345 13923 12403 13929
rect 12345 13889 12357 13923
rect 12391 13889 12403 13923
rect 12345 13883 12403 13889
rect 9122 13852 9128 13864
rect 8864 13824 9128 13852
rect 8573 13815 8631 13821
rect 9122 13812 9128 13824
rect 9180 13812 9186 13864
rect 9214 13812 9220 13864
rect 9272 13852 9278 13864
rect 9582 13852 9588 13864
rect 9272 13824 9588 13852
rect 9272 13816 9309 13824
rect 9272 13812 9278 13816
rect 9582 13812 9588 13824
rect 9640 13812 9646 13864
rect 10962 13812 10968 13864
rect 11020 13852 11026 13864
rect 11606 13852 11612 13864
rect 11020 13824 11612 13852
rect 11020 13812 11026 13824
rect 11606 13812 11612 13824
rect 11664 13812 11670 13864
rect 11698 13812 11704 13864
rect 11756 13852 11762 13864
rect 12360 13852 12388 13883
rect 12434 13880 12440 13932
rect 12492 13920 12498 13932
rect 12621 13923 12679 13929
rect 12621 13920 12633 13923
rect 12492 13892 12633 13920
rect 12492 13880 12498 13892
rect 12621 13889 12633 13892
rect 12667 13920 12679 13923
rect 12710 13920 12716 13932
rect 12667 13892 12716 13920
rect 12667 13889 12679 13892
rect 12621 13883 12679 13889
rect 12710 13880 12716 13892
rect 12768 13880 12774 13932
rect 13004 13929 13032 13960
rect 13906 13948 13912 14000
rect 13964 13988 13970 14000
rect 18417 13991 18475 13997
rect 18417 13988 18429 13991
rect 13964 13960 18429 13988
rect 13964 13948 13970 13960
rect 18417 13957 18429 13960
rect 18463 13957 18475 13991
rect 18417 13951 18475 13957
rect 12989 13923 13047 13929
rect 12989 13889 13001 13923
rect 13035 13920 13047 13923
rect 13170 13920 13176 13932
rect 13035 13892 13176 13920
rect 13035 13889 13047 13892
rect 12989 13883 13047 13889
rect 13170 13880 13176 13892
rect 13228 13880 13234 13932
rect 15746 13880 15752 13932
rect 15804 13920 15810 13932
rect 18049 13923 18107 13929
rect 18049 13920 18061 13923
rect 15804 13892 18061 13920
rect 15804 13880 15810 13892
rect 18049 13889 18061 13892
rect 18095 13889 18107 13923
rect 18049 13883 18107 13889
rect 18230 13880 18236 13932
rect 18288 13920 18294 13932
rect 19334 13920 19340 13932
rect 18288 13892 19340 13920
rect 18288 13880 18294 13892
rect 19334 13880 19340 13892
rect 19392 13880 19398 13932
rect 11756 13824 12388 13852
rect 11756 13812 11762 13824
rect 13722 13812 13728 13864
rect 13780 13852 13786 13864
rect 16574 13852 16580 13864
rect 13780 13824 16580 13852
rect 13780 13812 13786 13824
rect 16574 13812 16580 13824
rect 16632 13812 16638 13864
rect 9217 13807 9275 13812
rect 5040 13756 6684 13784
rect 5040 13744 5046 13756
rect 6730 13744 6736 13796
rect 6788 13784 6794 13796
rect 14550 13784 14556 13796
rect 6788 13756 9168 13784
rect 6788 13744 6794 13756
rect 3237 13719 3295 13725
rect 3237 13685 3249 13719
rect 3283 13716 3295 13719
rect 3602 13716 3608 13728
rect 3283 13688 3608 13716
rect 3283 13685 3295 13688
rect 3237 13679 3295 13685
rect 3602 13676 3608 13688
rect 3660 13676 3666 13728
rect 3970 13676 3976 13728
rect 4028 13716 4034 13728
rect 5077 13719 5135 13725
rect 5077 13716 5089 13719
rect 4028 13688 5089 13716
rect 4028 13676 4034 13688
rect 5077 13685 5089 13688
rect 5123 13685 5135 13719
rect 5077 13679 5135 13685
rect 5166 13676 5172 13728
rect 5224 13716 5230 13728
rect 5261 13719 5319 13725
rect 5261 13716 5273 13719
rect 5224 13688 5273 13716
rect 5224 13676 5230 13688
rect 5261 13685 5273 13688
rect 5307 13685 5319 13719
rect 5261 13679 5319 13685
rect 5718 13676 5724 13728
rect 5776 13676 5782 13728
rect 6270 13676 6276 13728
rect 6328 13716 6334 13728
rect 6822 13716 6828 13728
rect 6328 13688 6828 13716
rect 6328 13676 6334 13688
rect 6822 13676 6828 13688
rect 6880 13676 6886 13728
rect 7193 13719 7251 13725
rect 7193 13685 7205 13719
rect 7239 13716 7251 13719
rect 7558 13716 7564 13728
rect 7239 13688 7564 13716
rect 7239 13685 7251 13688
rect 7193 13679 7251 13685
rect 7558 13676 7564 13688
rect 7616 13716 7622 13728
rect 7926 13716 7932 13728
rect 7616 13688 7932 13716
rect 7616 13676 7622 13688
rect 7926 13676 7932 13688
rect 7984 13676 7990 13728
rect 8478 13676 8484 13728
rect 8536 13716 8542 13728
rect 9033 13719 9091 13725
rect 9033 13716 9045 13719
rect 8536 13688 9045 13716
rect 8536 13676 8542 13688
rect 9033 13685 9045 13688
rect 9079 13685 9091 13719
rect 9140 13716 9168 13756
rect 10336 13756 14556 13784
rect 10336 13716 10364 13756
rect 14550 13744 14556 13756
rect 14608 13744 14614 13796
rect 9140 13688 10364 13716
rect 9033 13679 9091 13685
rect 10410 13676 10416 13728
rect 10468 13716 10474 13728
rect 11422 13716 11428 13728
rect 10468 13688 11428 13716
rect 10468 13676 10474 13688
rect 11422 13676 11428 13688
rect 11480 13676 11486 13728
rect 12250 13676 12256 13728
rect 12308 13716 12314 13728
rect 12434 13716 12440 13728
rect 12308 13688 12440 13716
rect 12308 13676 12314 13688
rect 12434 13676 12440 13688
rect 12492 13676 12498 13728
rect 12526 13676 12532 13728
rect 12584 13716 12590 13728
rect 12621 13719 12679 13725
rect 12621 13716 12633 13719
rect 12584 13688 12633 13716
rect 12584 13676 12590 13688
rect 12621 13685 12633 13688
rect 12667 13685 12679 13719
rect 12621 13679 12679 13685
rect 12710 13676 12716 13728
rect 12768 13716 12774 13728
rect 13446 13716 13452 13728
rect 12768 13688 13452 13716
rect 12768 13676 12774 13688
rect 13446 13676 13452 13688
rect 13504 13676 13510 13728
rect 14918 13676 14924 13728
rect 14976 13716 14982 13728
rect 17126 13716 17132 13728
rect 14976 13688 17132 13716
rect 14976 13676 14982 13688
rect 17126 13676 17132 13688
rect 17184 13676 17190 13728
rect 1104 13626 18860 13648
rect 1104 13574 1950 13626
rect 2002 13574 2014 13626
rect 2066 13574 2078 13626
rect 2130 13574 2142 13626
rect 2194 13574 2206 13626
rect 2258 13574 6950 13626
rect 7002 13574 7014 13626
rect 7066 13574 7078 13626
rect 7130 13574 7142 13626
rect 7194 13574 7206 13626
rect 7258 13574 11950 13626
rect 12002 13574 12014 13626
rect 12066 13574 12078 13626
rect 12130 13574 12142 13626
rect 12194 13574 12206 13626
rect 12258 13574 16950 13626
rect 17002 13574 17014 13626
rect 17066 13574 17078 13626
rect 17130 13574 17142 13626
rect 17194 13574 17206 13626
rect 17258 13574 18860 13626
rect 1104 13552 18860 13574
rect 2222 13472 2228 13524
rect 2280 13512 2286 13524
rect 2280 13484 2774 13512
rect 2280 13472 2286 13484
rect 2746 13444 2774 13484
rect 3142 13472 3148 13524
rect 3200 13472 3206 13524
rect 4706 13472 4712 13524
rect 4764 13512 4770 13524
rect 4982 13512 4988 13524
rect 4764 13484 4988 13512
rect 4764 13472 4770 13484
rect 4982 13472 4988 13484
rect 5040 13472 5046 13524
rect 5169 13515 5227 13521
rect 5169 13481 5181 13515
rect 5215 13512 5227 13515
rect 5350 13512 5356 13524
rect 5215 13484 5356 13512
rect 5215 13481 5227 13484
rect 5169 13475 5227 13481
rect 5350 13472 5356 13484
rect 5408 13472 5414 13524
rect 5442 13472 5448 13524
rect 5500 13512 5506 13524
rect 9030 13512 9036 13524
rect 5500 13484 9036 13512
rect 5500 13472 5506 13484
rect 9030 13472 9036 13484
rect 9088 13472 9094 13524
rect 9490 13472 9496 13524
rect 9548 13472 9554 13524
rect 10042 13472 10048 13524
rect 10100 13512 10106 13524
rect 17218 13512 17224 13524
rect 10100 13484 17224 13512
rect 10100 13472 10106 13484
rect 17218 13472 17224 13484
rect 17276 13472 17282 13524
rect 18414 13472 18420 13524
rect 18472 13472 18478 13524
rect 6730 13444 6736 13456
rect 2746 13416 6736 13444
rect 6730 13404 6736 13416
rect 6788 13404 6794 13456
rect 8202 13444 8208 13456
rect 7024 13416 8208 13444
rect 934 13336 940 13388
rect 992 13376 998 13388
rect 5166 13376 5172 13388
rect 992 13348 5172 13376
rect 992 13336 998 13348
rect 5166 13336 5172 13348
rect 5224 13336 5230 13388
rect 5442 13336 5448 13388
rect 5500 13376 5506 13388
rect 5721 13379 5779 13385
rect 5721 13376 5733 13379
rect 5500 13348 5733 13376
rect 5500 13336 5506 13348
rect 5721 13345 5733 13348
rect 5767 13345 5779 13379
rect 5721 13339 5779 13345
rect 6086 13336 6092 13388
rect 6144 13336 6150 13388
rect 6454 13336 6460 13388
rect 6512 13376 6518 13388
rect 6914 13376 6920 13388
rect 6512 13348 6920 13376
rect 6512 13336 6518 13348
rect 6914 13336 6920 13348
rect 6972 13336 6978 13388
rect 2314 13268 2320 13320
rect 2372 13268 2378 13320
rect 2498 13268 2504 13320
rect 2556 13268 2562 13320
rect 2590 13268 2596 13320
rect 2648 13268 2654 13320
rect 2866 13268 2872 13320
rect 2924 13268 2930 13320
rect 2958 13268 2964 13320
rect 3016 13268 3022 13320
rect 3053 13311 3111 13317
rect 3053 13277 3065 13311
rect 3099 13308 3111 13311
rect 3142 13308 3148 13320
rect 3099 13280 3148 13308
rect 3099 13277 3111 13280
rect 3053 13271 3111 13277
rect 3142 13268 3148 13280
rect 3200 13268 3206 13320
rect 3237 13311 3295 13317
rect 3237 13277 3249 13311
rect 3283 13308 3295 13311
rect 4062 13308 4068 13320
rect 3283 13280 4068 13308
rect 3283 13277 3295 13280
rect 3237 13271 3295 13277
rect 4062 13268 4068 13280
rect 4120 13268 4126 13320
rect 4522 13268 4528 13320
rect 4580 13308 4586 13320
rect 5261 13311 5319 13317
rect 5261 13308 5273 13311
rect 4580 13280 5273 13308
rect 4580 13268 4586 13280
rect 5261 13277 5273 13280
rect 5307 13277 5319 13311
rect 5261 13271 5319 13277
rect 5997 13311 6055 13317
rect 5997 13277 6009 13311
rect 6043 13308 6055 13311
rect 6104 13308 6132 13336
rect 6043 13280 6132 13308
rect 6043 13277 6055 13280
rect 5997 13271 6055 13277
rect 6270 13268 6276 13320
rect 6328 13268 6334 13320
rect 7024 13317 7052 13416
rect 8202 13404 8208 13416
rect 8260 13404 8266 13456
rect 10226 13404 10232 13456
rect 10284 13444 10290 13456
rect 11054 13444 11060 13456
rect 10284 13416 11060 13444
rect 10284 13404 10290 13416
rect 11054 13404 11060 13416
rect 11112 13444 11118 13456
rect 12621 13447 12679 13453
rect 11112 13416 12572 13444
rect 11112 13404 11118 13416
rect 7101 13379 7159 13385
rect 7101 13345 7113 13379
rect 7147 13376 7159 13379
rect 7282 13376 7288 13388
rect 7147 13348 7288 13376
rect 7147 13345 7159 13348
rect 7101 13339 7159 13345
rect 7282 13336 7288 13348
rect 7340 13336 7346 13388
rect 7561 13379 7619 13385
rect 7561 13345 7573 13379
rect 7607 13376 7619 13379
rect 8110 13376 8116 13388
rect 7607 13348 8116 13376
rect 7607 13345 7619 13348
rect 7561 13339 7619 13345
rect 8110 13336 8116 13348
rect 8168 13376 8174 13388
rect 9306 13376 9312 13388
rect 8168 13348 9312 13376
rect 8168 13336 8174 13348
rect 9306 13336 9312 13348
rect 9364 13336 9370 13388
rect 9858 13376 9864 13388
rect 9692 13348 9864 13376
rect 7009 13311 7067 13317
rect 7009 13277 7021 13311
rect 7055 13277 7067 13311
rect 7009 13271 7067 13277
rect 7377 13311 7435 13317
rect 7377 13277 7389 13311
rect 7423 13308 7435 13311
rect 7926 13308 7932 13320
rect 7423 13280 7932 13308
rect 7423 13277 7435 13280
rect 7377 13271 7435 13277
rect 2332 13240 2360 13268
rect 2685 13243 2743 13249
rect 2685 13240 2697 13243
rect 2332 13212 2697 13240
rect 2685 13209 2697 13212
rect 2731 13209 2743 13243
rect 2685 13203 2743 13209
rect 1762 13132 1768 13184
rect 1820 13172 1826 13184
rect 2317 13175 2375 13181
rect 2317 13172 2329 13175
rect 1820 13144 2329 13172
rect 1820 13132 1826 13144
rect 2317 13141 2329 13144
rect 2363 13141 2375 13175
rect 2700 13172 2728 13203
rect 3786 13200 3792 13252
rect 3844 13240 3850 13252
rect 4246 13240 4252 13252
rect 3844 13212 4252 13240
rect 3844 13200 3850 13212
rect 4246 13200 4252 13212
rect 4304 13240 4310 13252
rect 5350 13240 5356 13252
rect 4304 13212 5356 13240
rect 4304 13200 4310 13212
rect 5350 13200 5356 13212
rect 5408 13200 5414 13252
rect 6086 13200 6092 13252
rect 6144 13240 6150 13252
rect 7392 13240 7420 13271
rect 7926 13268 7932 13280
rect 7984 13268 7990 13320
rect 8294 13268 8300 13320
rect 8352 13308 8358 13320
rect 9692 13317 9720 13348
rect 9858 13336 9864 13348
rect 9916 13336 9922 13388
rect 10870 13376 10876 13388
rect 10244 13348 10876 13376
rect 9677 13311 9735 13317
rect 9677 13308 9689 13311
rect 8352 13280 9689 13308
rect 8352 13268 8358 13280
rect 9677 13277 9689 13280
rect 9723 13277 9735 13311
rect 9677 13271 9735 13277
rect 9953 13311 10011 13317
rect 9953 13277 9965 13311
rect 9999 13308 10011 13311
rect 10244 13308 10272 13348
rect 10870 13336 10876 13348
rect 10928 13336 10934 13388
rect 11149 13379 11207 13385
rect 11149 13345 11161 13379
rect 11195 13376 11207 13379
rect 11882 13376 11888 13388
rect 11195 13348 11888 13376
rect 11195 13345 11207 13348
rect 11149 13339 11207 13345
rect 11882 13336 11888 13348
rect 11940 13336 11946 13388
rect 11974 13336 11980 13388
rect 12032 13376 12038 13388
rect 12434 13376 12440 13388
rect 12032 13348 12440 13376
rect 12032 13336 12038 13348
rect 12434 13336 12440 13348
rect 12492 13336 12498 13388
rect 12544 13376 12572 13416
rect 12621 13413 12633 13447
rect 12667 13444 12679 13447
rect 19426 13444 19432 13456
rect 12667 13416 19432 13444
rect 12667 13413 12679 13416
rect 12621 13407 12679 13413
rect 19426 13404 19432 13416
rect 19484 13404 19490 13456
rect 13998 13376 14004 13388
rect 12544 13348 14004 13376
rect 13998 13336 14004 13348
rect 14056 13336 14062 13388
rect 9999 13280 10272 13308
rect 9999 13277 10011 13280
rect 9953 13271 10011 13277
rect 11238 13268 11244 13320
rect 11296 13268 11302 13320
rect 12618 13268 12624 13320
rect 12676 13268 12682 13320
rect 12805 13311 12863 13317
rect 12805 13277 12817 13311
rect 12851 13277 12863 13311
rect 12805 13271 12863 13277
rect 12897 13311 12955 13317
rect 12897 13277 12909 13311
rect 12943 13308 12955 13311
rect 13078 13308 13084 13320
rect 12943 13280 13084 13308
rect 12943 13277 12955 13280
rect 12897 13271 12955 13277
rect 6144 13212 7420 13240
rect 8021 13243 8079 13249
rect 6144 13200 6150 13212
rect 8021 13209 8033 13243
rect 8067 13240 8079 13243
rect 8202 13240 8208 13252
rect 8067 13212 8208 13240
rect 8067 13209 8079 13212
rect 8021 13203 8079 13209
rect 8202 13200 8208 13212
rect 8260 13200 8266 13252
rect 9769 13243 9827 13249
rect 9769 13209 9781 13243
rect 9815 13240 9827 13243
rect 9858 13240 9864 13252
rect 9815 13212 9864 13240
rect 9815 13209 9827 13212
rect 9769 13203 9827 13209
rect 9858 13200 9864 13212
rect 9916 13200 9922 13252
rect 11790 13240 11796 13252
rect 11440 13212 11796 13240
rect 7006 13172 7012 13184
rect 2700 13144 7012 13172
rect 2317 13135 2375 13141
rect 7006 13132 7012 13144
rect 7064 13172 7070 13184
rect 11440 13172 11468 13212
rect 11790 13200 11796 13212
rect 11848 13240 11854 13252
rect 12820 13240 12848 13271
rect 13078 13268 13084 13280
rect 13136 13268 13142 13320
rect 13262 13268 13268 13320
rect 13320 13308 13326 13320
rect 13630 13308 13636 13320
rect 13320 13280 13636 13308
rect 13320 13268 13326 13280
rect 13630 13268 13636 13280
rect 13688 13268 13694 13320
rect 14642 13268 14648 13320
rect 14700 13308 14706 13320
rect 15105 13311 15163 13317
rect 15105 13308 15117 13311
rect 14700 13280 15117 13308
rect 14700 13268 14706 13280
rect 15105 13277 15117 13280
rect 15151 13277 15163 13311
rect 15105 13271 15163 13277
rect 15194 13268 15200 13320
rect 15252 13308 15258 13320
rect 15289 13311 15347 13317
rect 15289 13308 15301 13311
rect 15252 13280 15301 13308
rect 15252 13268 15258 13280
rect 15289 13277 15301 13280
rect 15335 13277 15347 13311
rect 15289 13271 15347 13277
rect 15470 13268 15476 13320
rect 15528 13268 15534 13320
rect 16666 13268 16672 13320
rect 16724 13308 16730 13320
rect 18049 13311 18107 13317
rect 16724 13280 17434 13308
rect 16724 13268 16730 13280
rect 18049 13277 18061 13311
rect 18095 13277 18107 13311
rect 18049 13271 18107 13277
rect 11848 13212 12848 13240
rect 11848 13200 11854 13212
rect 16850 13200 16856 13252
rect 16908 13240 16914 13252
rect 17037 13243 17095 13249
rect 17037 13240 17049 13243
rect 16908 13212 17049 13240
rect 16908 13200 16914 13212
rect 17037 13209 17049 13212
rect 17083 13209 17095 13243
rect 17037 13203 17095 13209
rect 17494 13200 17500 13252
rect 17552 13240 17558 13252
rect 18064 13240 18092 13271
rect 18230 13268 18236 13320
rect 18288 13268 18294 13320
rect 17552 13212 18092 13240
rect 17552 13200 17558 13212
rect 7064 13144 11468 13172
rect 7064 13132 7070 13144
rect 11606 13132 11612 13184
rect 11664 13132 11670 13184
rect 11698 13132 11704 13184
rect 11756 13172 11762 13184
rect 15838 13172 15844 13184
rect 11756 13144 15844 13172
rect 11756 13132 11762 13144
rect 15838 13132 15844 13144
rect 15896 13132 15902 13184
rect 1104 13082 18860 13104
rect 1104 13030 2610 13082
rect 2662 13030 2674 13082
rect 2726 13030 2738 13082
rect 2790 13030 2802 13082
rect 2854 13030 2866 13082
rect 2918 13030 7610 13082
rect 7662 13030 7674 13082
rect 7726 13030 7738 13082
rect 7790 13030 7802 13082
rect 7854 13030 7866 13082
rect 7918 13030 12610 13082
rect 12662 13030 12674 13082
rect 12726 13030 12738 13082
rect 12790 13030 12802 13082
rect 12854 13030 12866 13082
rect 12918 13030 17610 13082
rect 17662 13030 17674 13082
rect 17726 13030 17738 13082
rect 17790 13030 17802 13082
rect 17854 13030 17866 13082
rect 17918 13030 18860 13082
rect 1104 13008 18860 13030
rect 2314 12928 2320 12980
rect 2372 12968 2378 12980
rect 2682 12968 2688 12980
rect 2372 12940 2688 12968
rect 2372 12928 2378 12940
rect 2682 12928 2688 12940
rect 2740 12928 2746 12980
rect 2958 12928 2964 12980
rect 3016 12968 3022 12980
rect 6457 12971 6515 12977
rect 6457 12968 6469 12971
rect 3016 12940 6469 12968
rect 3016 12928 3022 12940
rect 6457 12937 6469 12940
rect 6503 12937 6515 12971
rect 6457 12931 6515 12937
rect 7374 12928 7380 12980
rect 7432 12968 7438 12980
rect 7561 12971 7619 12977
rect 7561 12968 7573 12971
rect 7432 12940 7573 12968
rect 7432 12928 7438 12940
rect 7561 12937 7573 12940
rect 7607 12937 7619 12971
rect 7561 12931 7619 12937
rect 7650 12928 7656 12980
rect 7708 12968 7714 12980
rect 7745 12971 7803 12977
rect 7745 12968 7757 12971
rect 7708 12940 7757 12968
rect 7708 12928 7714 12940
rect 7745 12937 7757 12940
rect 7791 12937 7803 12971
rect 7745 12931 7803 12937
rect 9214 12928 9220 12980
rect 9272 12968 9278 12980
rect 11514 12968 11520 12980
rect 9272 12940 11520 12968
rect 9272 12928 9278 12940
rect 11514 12928 11520 12940
rect 11572 12928 11578 12980
rect 11882 12928 11888 12980
rect 11940 12968 11946 12980
rect 12805 12971 12863 12977
rect 12805 12968 12817 12971
rect 11940 12940 12817 12968
rect 11940 12928 11946 12940
rect 12805 12937 12817 12940
rect 12851 12968 12863 12971
rect 15010 12968 15016 12980
rect 12851 12940 15016 12968
rect 12851 12937 12863 12940
rect 12805 12931 12863 12937
rect 15010 12928 15016 12940
rect 15068 12928 15074 12980
rect 15286 12928 15292 12980
rect 15344 12968 15350 12980
rect 15470 12968 15476 12980
rect 15344 12940 15476 12968
rect 15344 12928 15350 12940
rect 15470 12928 15476 12940
rect 15528 12928 15534 12980
rect 16022 12928 16028 12980
rect 16080 12968 16086 12980
rect 18046 12968 18052 12980
rect 16080 12940 18052 12968
rect 16080 12928 16086 12940
rect 18046 12928 18052 12940
rect 18104 12928 18110 12980
rect 1946 12860 1952 12912
rect 2004 12900 2010 12912
rect 2222 12900 2228 12912
rect 2004 12872 2228 12900
rect 2004 12860 2010 12872
rect 2222 12860 2228 12872
rect 2280 12900 2286 12912
rect 3329 12903 3387 12909
rect 3329 12900 3341 12903
rect 2280 12872 3341 12900
rect 2280 12860 2286 12872
rect 3329 12869 3341 12872
rect 3375 12869 3387 12903
rect 3329 12863 3387 12869
rect 3421 12903 3479 12909
rect 3421 12869 3433 12903
rect 3467 12900 3479 12903
rect 3510 12900 3516 12912
rect 3467 12872 3516 12900
rect 3467 12869 3479 12872
rect 3421 12863 3479 12869
rect 3510 12860 3516 12872
rect 3568 12860 3574 12912
rect 4157 12903 4215 12909
rect 4157 12869 4169 12903
rect 4203 12900 4215 12903
rect 4706 12900 4712 12912
rect 4203 12872 4712 12900
rect 4203 12869 4215 12872
rect 4157 12863 4215 12869
rect 4706 12860 4712 12872
rect 4764 12860 4770 12912
rect 4982 12860 4988 12912
rect 5040 12860 5046 12912
rect 9861 12903 9919 12909
rect 9861 12900 9873 12903
rect 5184 12872 9873 12900
rect 2593 12835 2651 12841
rect 2593 12801 2605 12835
rect 2639 12832 2651 12835
rect 2774 12832 2780 12844
rect 2639 12804 2780 12832
rect 2639 12801 2651 12804
rect 2593 12795 2651 12801
rect 2774 12792 2780 12804
rect 2832 12792 2838 12844
rect 3050 12792 3056 12844
rect 3108 12792 3114 12844
rect 3234 12792 3240 12844
rect 3292 12792 3298 12844
rect 3697 12835 3755 12841
rect 3697 12801 3709 12835
rect 3743 12801 3755 12835
rect 3697 12795 3755 12801
rect 474 12724 480 12776
rect 532 12764 538 12776
rect 1854 12764 1860 12776
rect 532 12736 1860 12764
rect 532 12724 538 12736
rect 1854 12724 1860 12736
rect 1912 12724 1918 12776
rect 2498 12724 2504 12776
rect 2556 12724 2562 12776
rect 2958 12724 2964 12776
rect 3016 12724 3022 12776
rect 3068 12764 3096 12792
rect 3712 12764 3740 12795
rect 4614 12792 4620 12844
rect 4672 12792 4678 12844
rect 5184 12841 5212 12872
rect 9861 12869 9873 12872
rect 9907 12900 9919 12903
rect 10410 12900 10416 12912
rect 9907 12872 10416 12900
rect 9907 12869 9919 12872
rect 9861 12863 9919 12869
rect 10410 12860 10416 12872
rect 10468 12860 10474 12912
rect 13078 12900 13084 12912
rect 10704 12872 13084 12900
rect 5169 12835 5227 12841
rect 5169 12801 5181 12835
rect 5215 12801 5227 12835
rect 5169 12795 5227 12801
rect 5350 12792 5356 12844
rect 5408 12792 5414 12844
rect 5442 12792 5448 12844
rect 5500 12792 5506 12844
rect 5626 12792 5632 12844
rect 5684 12832 5690 12844
rect 6546 12832 6552 12844
rect 5684 12804 6552 12832
rect 5684 12792 5690 12804
rect 6546 12792 6552 12804
rect 6604 12832 6610 12844
rect 6641 12835 6699 12841
rect 6641 12832 6653 12835
rect 6604 12804 6653 12832
rect 6604 12792 6610 12804
rect 6641 12801 6653 12804
rect 6687 12801 6699 12835
rect 6641 12795 6699 12801
rect 6730 12792 6736 12844
rect 6788 12792 6794 12844
rect 7006 12792 7012 12844
rect 7064 12792 7070 12844
rect 7558 12792 7564 12844
rect 7616 12832 7622 12844
rect 7616 12804 7661 12832
rect 7616 12792 7622 12804
rect 7742 12792 7748 12844
rect 7800 12832 7806 12844
rect 8386 12832 8392 12844
rect 7800 12804 8392 12832
rect 7800 12792 7806 12804
rect 8386 12792 8392 12804
rect 8444 12792 8450 12844
rect 9306 12792 9312 12844
rect 9364 12832 9370 12844
rect 9364 12804 9904 12832
rect 9364 12792 9370 12804
rect 3068 12736 3740 12764
rect 3712 12696 3740 12736
rect 4525 12767 4583 12773
rect 4525 12733 4537 12767
rect 4571 12733 4583 12767
rect 4525 12727 4583 12733
rect 7101 12767 7159 12773
rect 7101 12733 7113 12767
rect 7147 12764 7159 12767
rect 8294 12764 8300 12776
rect 7147 12736 8300 12764
rect 7147 12733 7159 12736
rect 7101 12727 7159 12733
rect 4540 12696 4568 12727
rect 8294 12724 8300 12736
rect 8352 12724 8358 12776
rect 9030 12724 9036 12776
rect 9088 12764 9094 12776
rect 9766 12764 9772 12776
rect 9088 12736 9772 12764
rect 9088 12724 9094 12736
rect 9766 12724 9772 12736
rect 9824 12724 9830 12776
rect 9876 12764 9904 12804
rect 10042 12792 10048 12844
rect 10100 12792 10106 12844
rect 10704 12832 10732 12872
rect 13078 12860 13084 12872
rect 13136 12860 13142 12912
rect 13262 12860 13268 12912
rect 13320 12900 13326 12912
rect 13320 12872 16160 12900
rect 13320 12860 13326 12872
rect 10428 12804 10732 12832
rect 10781 12835 10839 12841
rect 10428 12776 10456 12804
rect 10781 12801 10793 12835
rect 10827 12822 10839 12835
rect 10870 12822 10876 12844
rect 10827 12801 10876 12822
rect 10781 12795 10876 12801
rect 10796 12794 10876 12795
rect 10870 12792 10876 12794
rect 10928 12792 10934 12844
rect 10962 12792 10968 12844
rect 11020 12792 11026 12844
rect 11057 12835 11115 12841
rect 11057 12801 11069 12835
rect 11103 12832 11115 12835
rect 11238 12832 11244 12844
rect 11103 12804 11244 12832
rect 11103 12801 11115 12804
rect 11057 12795 11115 12801
rect 11238 12792 11244 12804
rect 11296 12792 11302 12844
rect 11330 12792 11336 12844
rect 11388 12832 11394 12844
rect 11517 12835 11575 12841
rect 11517 12832 11529 12835
rect 11388 12804 11529 12832
rect 11388 12792 11394 12804
rect 11517 12801 11529 12804
rect 11563 12801 11575 12835
rect 11517 12795 11575 12801
rect 11974 12792 11980 12844
rect 12032 12792 12038 12844
rect 12066 12792 12072 12844
rect 12124 12832 12130 12844
rect 12345 12835 12403 12841
rect 12345 12832 12357 12835
rect 12124 12804 12357 12832
rect 12124 12792 12130 12804
rect 12345 12801 12357 12804
rect 12391 12801 12403 12835
rect 12345 12795 12403 12801
rect 10137 12767 10195 12773
rect 10137 12764 10149 12767
rect 9876 12736 10149 12764
rect 10137 12733 10149 12736
rect 10183 12764 10195 12767
rect 10410 12764 10416 12776
rect 10183 12736 10416 12764
rect 10183 12733 10195 12736
rect 10137 12727 10195 12733
rect 10410 12724 10416 12736
rect 10468 12724 10474 12776
rect 10505 12767 10563 12773
rect 10505 12733 10517 12767
rect 10551 12764 10563 12767
rect 11698 12764 11704 12776
rect 10551 12736 11704 12764
rect 10551 12733 10563 12736
rect 10505 12727 10563 12733
rect 4614 12696 4620 12708
rect 3712 12668 4479 12696
rect 4540 12668 4620 12696
rect 2317 12631 2375 12637
rect 2317 12597 2329 12631
rect 2363 12628 2375 12631
rect 3234 12628 3240 12640
rect 2363 12600 3240 12628
rect 2363 12597 2375 12600
rect 2317 12591 2375 12597
rect 3234 12588 3240 12600
rect 3292 12588 3298 12640
rect 3602 12588 3608 12640
rect 3660 12588 3666 12640
rect 3878 12588 3884 12640
rect 3936 12588 3942 12640
rect 4451 12628 4479 12668
rect 4614 12656 4620 12668
rect 4672 12656 4678 12708
rect 4801 12699 4859 12705
rect 4801 12665 4813 12699
rect 4847 12696 4859 12699
rect 7558 12696 7564 12708
rect 4847 12668 7564 12696
rect 4847 12665 4859 12668
rect 4801 12659 4859 12665
rect 7558 12656 7564 12668
rect 7616 12656 7622 12708
rect 7742 12656 7748 12708
rect 7800 12696 7806 12708
rect 9582 12696 9588 12708
rect 7800 12668 9588 12696
rect 7800 12656 7806 12668
rect 9582 12656 9588 12668
rect 9640 12656 9646 12708
rect 9950 12656 9956 12708
rect 10008 12696 10014 12708
rect 10520 12696 10548 12727
rect 11698 12724 11704 12736
rect 11756 12724 11762 12776
rect 11790 12724 11796 12776
rect 11848 12764 11854 12776
rect 11885 12767 11943 12773
rect 11885 12764 11897 12767
rect 11848 12736 11897 12764
rect 11848 12724 11854 12736
rect 11885 12733 11897 12736
rect 11931 12733 11943 12767
rect 11885 12727 11943 12733
rect 12161 12767 12219 12773
rect 12161 12733 12173 12767
rect 12207 12764 12219 12767
rect 12250 12764 12256 12776
rect 12207 12736 12256 12764
rect 12207 12733 12219 12736
rect 12161 12727 12219 12733
rect 12250 12724 12256 12736
rect 12308 12724 12314 12776
rect 12360 12764 12388 12795
rect 12434 12792 12440 12844
rect 12492 12832 12498 12844
rect 12621 12835 12679 12841
rect 12621 12832 12633 12835
rect 12492 12804 12633 12832
rect 12492 12792 12498 12804
rect 12621 12801 12633 12804
rect 12667 12801 12679 12835
rect 12621 12795 12679 12801
rect 12894 12792 12900 12844
rect 12952 12832 12958 12844
rect 13446 12832 13452 12844
rect 12952 12804 13452 12832
rect 12952 12792 12958 12804
rect 13446 12792 13452 12804
rect 13504 12792 13510 12844
rect 14826 12792 14832 12844
rect 14884 12832 14890 12844
rect 15010 12832 15016 12844
rect 14884 12804 15016 12832
rect 14884 12792 14890 12804
rect 15010 12792 15016 12804
rect 15068 12792 15074 12844
rect 16022 12832 16028 12844
rect 15856 12804 16028 12832
rect 12710 12764 12716 12776
rect 12360 12736 12716 12764
rect 12710 12724 12716 12736
rect 12768 12724 12774 12776
rect 13906 12724 13912 12776
rect 13964 12764 13970 12776
rect 15856 12764 15884 12804
rect 16022 12792 16028 12804
rect 16080 12792 16086 12844
rect 16132 12841 16160 12872
rect 16298 12860 16304 12912
rect 16356 12900 16362 12912
rect 16356 12872 18092 12900
rect 16356 12860 16362 12872
rect 16117 12835 16175 12841
rect 16117 12801 16129 12835
rect 16163 12801 16175 12835
rect 16117 12795 16175 12801
rect 16209 12835 16267 12841
rect 16209 12801 16221 12835
rect 16255 12832 16267 12835
rect 16255 12804 16436 12832
rect 16255 12801 16267 12804
rect 16209 12795 16267 12801
rect 13964 12736 15884 12764
rect 13964 12724 13970 12736
rect 15930 12724 15936 12776
rect 15988 12764 15994 12776
rect 16301 12767 16359 12773
rect 16301 12764 16313 12767
rect 15988 12736 16313 12764
rect 15988 12724 15994 12736
rect 16301 12733 16313 12736
rect 16347 12733 16359 12767
rect 16301 12727 16359 12733
rect 10008 12668 10548 12696
rect 10008 12656 10014 12668
rect 10594 12656 10600 12708
rect 10652 12656 10658 12708
rect 12437 12699 12495 12705
rect 12437 12665 12449 12699
rect 12483 12665 12495 12699
rect 12437 12659 12495 12665
rect 12529 12699 12587 12705
rect 12529 12665 12541 12699
rect 12575 12696 12587 12699
rect 13170 12696 13176 12708
rect 12575 12668 13176 12696
rect 12575 12665 12587 12668
rect 12529 12659 12587 12665
rect 6730 12628 6736 12640
rect 4451 12600 6736 12628
rect 6730 12588 6736 12600
rect 6788 12588 6794 12640
rect 6822 12588 6828 12640
rect 6880 12628 6886 12640
rect 6917 12631 6975 12637
rect 6917 12628 6929 12631
rect 6880 12600 6929 12628
rect 6880 12588 6886 12600
rect 6917 12597 6929 12600
rect 6963 12597 6975 12631
rect 6917 12591 6975 12597
rect 7006 12588 7012 12640
rect 7064 12628 7070 12640
rect 7193 12631 7251 12637
rect 7193 12628 7205 12631
rect 7064 12600 7205 12628
rect 7064 12588 7070 12600
rect 7193 12597 7205 12600
rect 7239 12597 7251 12631
rect 7193 12591 7251 12597
rect 8386 12588 8392 12640
rect 8444 12628 8450 12640
rect 10502 12628 10508 12640
rect 8444 12600 10508 12628
rect 8444 12588 8450 12600
rect 10502 12588 10508 12600
rect 10560 12588 10566 12640
rect 10686 12588 10692 12640
rect 10744 12628 10750 12640
rect 11146 12628 11152 12640
rect 10744 12600 11152 12628
rect 10744 12588 10750 12600
rect 11146 12588 11152 12600
rect 11204 12588 11210 12640
rect 11238 12588 11244 12640
rect 11296 12628 11302 12640
rect 12452 12628 12480 12659
rect 13170 12656 13176 12668
rect 13228 12696 13234 12708
rect 13446 12696 13452 12708
rect 13228 12668 13452 12696
rect 13228 12656 13234 12668
rect 13446 12656 13452 12668
rect 13504 12696 13510 12708
rect 16408 12696 16436 12804
rect 17218 12792 17224 12844
rect 17276 12832 17282 12844
rect 17313 12835 17371 12841
rect 17313 12832 17325 12835
rect 17276 12804 17325 12832
rect 17276 12792 17282 12804
rect 17313 12801 17325 12804
rect 17359 12801 17371 12835
rect 17313 12795 17371 12801
rect 17328 12764 17356 12795
rect 17678 12792 17684 12844
rect 17736 12792 17742 12844
rect 18064 12841 18092 12872
rect 18322 12860 18328 12912
rect 18380 12900 18386 12912
rect 18417 12903 18475 12909
rect 18417 12900 18429 12903
rect 18380 12872 18429 12900
rect 18380 12860 18386 12872
rect 18417 12869 18429 12872
rect 18463 12869 18475 12903
rect 18417 12863 18475 12869
rect 18049 12835 18107 12841
rect 18049 12801 18061 12835
rect 18095 12801 18107 12835
rect 18049 12795 18107 12801
rect 18230 12764 18236 12776
rect 17328 12736 18236 12764
rect 18230 12724 18236 12736
rect 18288 12724 18294 12776
rect 13504 12668 16436 12696
rect 13504 12656 13510 12668
rect 11296 12600 12480 12628
rect 11296 12588 11302 12600
rect 12618 12588 12624 12640
rect 12676 12628 12682 12640
rect 13538 12628 13544 12640
rect 12676 12600 13544 12628
rect 12676 12588 12682 12600
rect 13538 12588 13544 12600
rect 13596 12588 13602 12640
rect 14182 12588 14188 12640
rect 14240 12628 14246 12640
rect 16485 12631 16543 12637
rect 16485 12628 16497 12631
rect 14240 12600 16497 12628
rect 14240 12588 14246 12600
rect 16485 12597 16497 12600
rect 16531 12597 16543 12631
rect 16485 12591 16543 12597
rect 17402 12588 17408 12640
rect 17460 12628 17466 12640
rect 18506 12628 18512 12640
rect 17460 12600 18512 12628
rect 17460 12588 17466 12600
rect 18506 12588 18512 12600
rect 18564 12588 18570 12640
rect 1104 12538 18860 12560
rect 1104 12486 1950 12538
rect 2002 12486 2014 12538
rect 2066 12486 2078 12538
rect 2130 12486 2142 12538
rect 2194 12486 2206 12538
rect 2258 12486 6950 12538
rect 7002 12486 7014 12538
rect 7066 12486 7078 12538
rect 7130 12486 7142 12538
rect 7194 12486 7206 12538
rect 7258 12486 11950 12538
rect 12002 12486 12014 12538
rect 12066 12486 12078 12538
rect 12130 12486 12142 12538
rect 12194 12486 12206 12538
rect 12258 12486 16950 12538
rect 17002 12486 17014 12538
rect 17066 12486 17078 12538
rect 17130 12486 17142 12538
rect 17194 12486 17206 12538
rect 17258 12486 18860 12538
rect 1104 12464 18860 12486
rect 2130 12384 2136 12436
rect 2188 12424 2194 12436
rect 3786 12424 3792 12436
rect 2188 12396 3792 12424
rect 2188 12384 2194 12396
rect 3786 12384 3792 12396
rect 3844 12384 3850 12436
rect 4154 12384 4160 12436
rect 4212 12424 4218 12436
rect 5626 12424 5632 12436
rect 4212 12396 5632 12424
rect 4212 12384 4218 12396
rect 5626 12384 5632 12396
rect 5684 12384 5690 12436
rect 5810 12384 5816 12436
rect 5868 12424 5874 12436
rect 7650 12424 7656 12436
rect 5868 12396 7656 12424
rect 5868 12384 5874 12396
rect 7650 12384 7656 12396
rect 7708 12384 7714 12436
rect 8202 12384 8208 12436
rect 8260 12424 8266 12436
rect 9030 12424 9036 12436
rect 8260 12396 9036 12424
rect 8260 12384 8266 12396
rect 9030 12384 9036 12396
rect 9088 12384 9094 12436
rect 9309 12427 9367 12433
rect 9309 12393 9321 12427
rect 9355 12424 9367 12427
rect 9766 12424 9772 12436
rect 9355 12396 9772 12424
rect 9355 12393 9367 12396
rect 9309 12387 9367 12393
rect 9766 12384 9772 12396
rect 9824 12384 9830 12436
rect 10134 12384 10140 12436
rect 10192 12424 10198 12436
rect 10689 12427 10747 12433
rect 10689 12424 10701 12427
rect 10192 12396 10701 12424
rect 10192 12384 10198 12396
rect 10689 12393 10701 12396
rect 10735 12393 10747 12427
rect 10689 12387 10747 12393
rect 12713 12427 12771 12433
rect 12713 12393 12725 12427
rect 12759 12424 12771 12427
rect 12986 12424 12992 12436
rect 12759 12396 12992 12424
rect 12759 12393 12771 12396
rect 12713 12387 12771 12393
rect 12986 12384 12992 12396
rect 13044 12384 13050 12436
rect 13538 12384 13544 12436
rect 13596 12424 13602 12436
rect 14826 12424 14832 12436
rect 13596 12396 14832 12424
rect 13596 12384 13602 12396
rect 14826 12384 14832 12396
rect 14884 12384 14890 12436
rect 15102 12384 15108 12436
rect 15160 12424 15166 12436
rect 16117 12427 16175 12433
rect 16117 12424 16129 12427
rect 15160 12396 16129 12424
rect 15160 12384 15166 12396
rect 16117 12393 16129 12396
rect 16163 12393 16175 12427
rect 16117 12387 16175 12393
rect 16206 12384 16212 12436
rect 16264 12424 16270 12436
rect 16853 12427 16911 12433
rect 16264 12396 16528 12424
rect 16264 12384 16270 12396
rect 16500 12368 16528 12396
rect 16853 12393 16865 12427
rect 16899 12424 16911 12427
rect 16899 12396 17448 12424
rect 16899 12393 16911 12396
rect 16853 12387 16911 12393
rect 4341 12359 4399 12365
rect 4341 12325 4353 12359
rect 4387 12356 4399 12359
rect 8110 12356 8116 12368
rect 4387 12328 8116 12356
rect 4387 12325 4399 12328
rect 4341 12319 4399 12325
rect 8110 12316 8116 12328
rect 8168 12316 8174 12368
rect 8938 12316 8944 12368
rect 8996 12356 9002 12368
rect 9674 12356 9680 12368
rect 8996 12328 9680 12356
rect 8996 12316 9002 12328
rect 9674 12316 9680 12328
rect 9732 12316 9738 12368
rect 10318 12316 10324 12368
rect 10376 12356 10382 12368
rect 11238 12356 11244 12368
rect 10376 12328 11244 12356
rect 10376 12316 10382 12328
rect 11238 12316 11244 12328
rect 11296 12316 11302 12368
rect 11330 12316 11336 12368
rect 11388 12356 11394 12368
rect 13265 12359 13323 12365
rect 13265 12356 13277 12359
rect 11388 12328 13277 12356
rect 11388 12316 11394 12328
rect 13265 12325 13277 12328
rect 13311 12325 13323 12359
rect 14642 12356 14648 12368
rect 13265 12319 13323 12325
rect 13556 12328 14648 12356
rect 13556 12300 13584 12328
rect 14642 12316 14648 12328
rect 14700 12316 14706 12368
rect 15746 12316 15752 12368
rect 15804 12356 15810 12368
rect 16393 12359 16451 12365
rect 16393 12356 16405 12359
rect 15804 12328 16405 12356
rect 15804 12316 15810 12328
rect 16393 12325 16405 12328
rect 16439 12325 16451 12359
rect 16393 12319 16451 12325
rect 16482 12316 16488 12368
rect 16540 12316 16546 12368
rect 17420 12356 17448 12396
rect 17494 12384 17500 12436
rect 17552 12424 17558 12436
rect 17865 12427 17923 12433
rect 17865 12424 17877 12427
rect 17552 12396 17877 12424
rect 17552 12384 17558 12396
rect 17865 12393 17877 12396
rect 17911 12393 17923 12427
rect 17865 12387 17923 12393
rect 18138 12356 18144 12368
rect 17420 12328 18144 12356
rect 18138 12316 18144 12328
rect 18196 12316 18202 12368
rect 1302 12248 1308 12300
rect 1360 12288 1366 12300
rect 3694 12288 3700 12300
rect 1360 12260 3700 12288
rect 1360 12248 1366 12260
rect 3694 12248 3700 12260
rect 3752 12288 3758 12300
rect 3789 12291 3847 12297
rect 3789 12288 3801 12291
rect 3752 12260 3801 12288
rect 3752 12248 3758 12260
rect 3789 12257 3801 12260
rect 3835 12257 3847 12291
rect 3789 12251 3847 12257
rect 5902 12248 5908 12300
rect 5960 12248 5966 12300
rect 5994 12248 6000 12300
rect 6052 12288 6058 12300
rect 7006 12288 7012 12300
rect 6052 12260 7012 12288
rect 6052 12248 6058 12260
rect 7006 12248 7012 12260
rect 7064 12248 7070 12300
rect 7282 12248 7288 12300
rect 7340 12288 7346 12300
rect 7340 12260 10824 12288
rect 7340 12248 7346 12260
rect 1394 12180 1400 12232
rect 1452 12220 1458 12232
rect 2409 12223 2467 12229
rect 2409 12220 2421 12223
rect 1452 12192 2421 12220
rect 1452 12180 1458 12192
rect 2409 12189 2421 12192
rect 2455 12189 2467 12223
rect 2409 12183 2467 12189
rect 3973 12223 4031 12229
rect 3973 12189 3985 12223
rect 4019 12189 4031 12223
rect 3973 12183 4031 12189
rect 2682 12112 2688 12164
rect 2740 12152 2746 12164
rect 2961 12155 3019 12161
rect 2961 12152 2973 12155
rect 2740 12124 2973 12152
rect 2740 12112 2746 12124
rect 2961 12121 2973 12124
rect 3007 12152 3019 12155
rect 3326 12152 3332 12164
rect 3007 12124 3332 12152
rect 3007 12121 3019 12124
rect 2961 12115 3019 12121
rect 3326 12112 3332 12124
rect 3384 12112 3390 12164
rect 3694 12112 3700 12164
rect 3752 12152 3758 12164
rect 3988 12152 4016 12183
rect 4246 12180 4252 12232
rect 4304 12220 4310 12232
rect 4430 12220 4436 12232
rect 4304 12192 4436 12220
rect 4304 12180 4310 12192
rect 4430 12180 4436 12192
rect 4488 12180 4494 12232
rect 4982 12180 4988 12232
rect 5040 12220 5046 12232
rect 5353 12223 5411 12229
rect 5353 12220 5365 12223
rect 5040 12192 5365 12220
rect 5040 12180 5046 12192
rect 5353 12189 5365 12192
rect 5399 12220 5411 12223
rect 5442 12220 5448 12232
rect 5399 12192 5448 12220
rect 5399 12189 5411 12192
rect 5353 12183 5411 12189
rect 5442 12180 5448 12192
rect 5500 12180 5506 12232
rect 6178 12180 6184 12232
rect 6236 12220 6242 12232
rect 6236 12216 6776 12220
rect 6932 12216 9168 12220
rect 6236 12192 9168 12216
rect 6236 12180 6242 12192
rect 6748 12188 6960 12192
rect 3752 12124 4016 12152
rect 4617 12155 4675 12161
rect 3752 12112 3758 12124
rect 4617 12121 4629 12155
rect 4663 12152 4675 12155
rect 5626 12152 5632 12164
rect 4663 12124 5632 12152
rect 4663 12121 4675 12124
rect 4617 12115 4675 12121
rect 5626 12112 5632 12124
rect 5684 12112 5690 12164
rect 6546 12112 6552 12164
rect 6604 12152 6610 12164
rect 7374 12152 7380 12164
rect 6604 12124 7380 12152
rect 6604 12112 6610 12124
rect 7374 12112 7380 12124
rect 7432 12152 7438 12164
rect 8754 12152 8760 12164
rect 7432 12124 8760 12152
rect 7432 12112 7438 12124
rect 8754 12112 8760 12124
rect 8812 12112 8818 12164
rect 9140 12152 9168 12192
rect 9214 12180 9220 12232
rect 9272 12180 9278 12232
rect 10226 12220 10232 12232
rect 9416 12192 10232 12220
rect 9306 12152 9312 12164
rect 9140 12124 9312 12152
rect 9306 12112 9312 12124
rect 9364 12112 9370 12164
rect 3510 12044 3516 12096
rect 3568 12084 3574 12096
rect 9416 12084 9444 12192
rect 10226 12180 10232 12192
rect 10284 12180 10290 12232
rect 10597 12223 10655 12229
rect 10597 12189 10609 12223
rect 10643 12220 10655 12223
rect 10686 12220 10692 12232
rect 10643 12192 10692 12220
rect 10643 12189 10655 12192
rect 10597 12183 10655 12189
rect 10686 12180 10692 12192
rect 10744 12180 10750 12232
rect 10796 12229 10824 12260
rect 11606 12248 11612 12300
rect 11664 12288 11670 12300
rect 12434 12288 12440 12300
rect 11664 12260 12440 12288
rect 11664 12248 11670 12260
rect 12434 12248 12440 12260
rect 12492 12248 12498 12300
rect 13078 12288 13084 12300
rect 12912 12260 13084 12288
rect 10781 12223 10839 12229
rect 10781 12189 10793 12223
rect 10827 12220 10839 12223
rect 12618 12220 12624 12232
rect 10827 12192 12624 12220
rect 10827 12189 10839 12192
rect 10781 12183 10839 12189
rect 12618 12180 12624 12192
rect 12676 12180 12682 12232
rect 12912 12229 12940 12260
rect 13078 12248 13084 12260
rect 13136 12248 13142 12300
rect 13538 12248 13544 12300
rect 13596 12248 13602 12300
rect 16942 12288 16948 12300
rect 13648 12260 16948 12288
rect 12897 12223 12955 12229
rect 12897 12189 12909 12223
rect 12943 12189 12955 12223
rect 12897 12183 12955 12189
rect 12986 12180 12992 12232
rect 13044 12180 13050 12232
rect 13170 12180 13176 12232
rect 13228 12180 13234 12232
rect 13449 12223 13507 12229
rect 13449 12189 13461 12223
rect 13495 12189 13507 12223
rect 13449 12183 13507 12189
rect 9582 12112 9588 12164
rect 9640 12152 9646 12164
rect 12345 12155 12403 12161
rect 12345 12152 12357 12155
rect 9640 12124 12357 12152
rect 9640 12112 9646 12124
rect 12345 12121 12357 12124
rect 12391 12121 12403 12155
rect 12345 12115 12403 12121
rect 12529 12155 12587 12161
rect 12529 12121 12541 12155
rect 12575 12152 12587 12155
rect 13464 12152 13492 12183
rect 13648 12152 13676 12260
rect 16942 12248 16948 12260
rect 17000 12248 17006 12300
rect 17402 12248 17408 12300
rect 17460 12248 17466 12300
rect 17512 12260 18552 12288
rect 14461 12223 14519 12229
rect 14461 12189 14473 12223
rect 14507 12189 14519 12223
rect 14461 12183 14519 12189
rect 14645 12223 14703 12229
rect 14645 12189 14657 12223
rect 14691 12220 14703 12223
rect 15378 12220 15384 12232
rect 14691 12192 15384 12220
rect 14691 12189 14703 12192
rect 14645 12183 14703 12189
rect 12575 12124 13676 12152
rect 12575 12121 12587 12124
rect 12529 12115 12587 12121
rect 13998 12112 14004 12164
rect 14056 12152 14062 12164
rect 14093 12155 14151 12161
rect 14093 12152 14105 12155
rect 14056 12124 14105 12152
rect 14056 12112 14062 12124
rect 14093 12121 14105 12124
rect 14139 12121 14151 12155
rect 14093 12115 14151 12121
rect 14185 12155 14243 12161
rect 14185 12121 14197 12155
rect 14231 12152 14243 12155
rect 14274 12152 14280 12164
rect 14231 12124 14280 12152
rect 14231 12121 14243 12124
rect 14185 12115 14243 12121
rect 3568 12056 9444 12084
rect 3568 12044 3574 12056
rect 9766 12044 9772 12096
rect 9824 12084 9830 12096
rect 10778 12084 10784 12096
rect 9824 12056 10784 12084
rect 9824 12044 9830 12056
rect 10778 12044 10784 12056
rect 10836 12044 10842 12096
rect 12250 12044 12256 12096
rect 12308 12084 12314 12096
rect 12710 12084 12716 12096
rect 12308 12056 12716 12084
rect 12308 12044 12314 12056
rect 12710 12044 12716 12056
rect 12768 12044 12774 12096
rect 13170 12044 13176 12096
rect 13228 12084 13234 12096
rect 13354 12084 13360 12096
rect 13228 12056 13360 12084
rect 13228 12044 13234 12056
rect 13354 12044 13360 12056
rect 13412 12044 13418 12096
rect 14108 12084 14136 12115
rect 14274 12112 14280 12124
rect 14332 12112 14338 12164
rect 14476 12152 14504 12183
rect 15378 12180 15384 12192
rect 15436 12180 15442 12232
rect 16298 12180 16304 12232
rect 16356 12180 16362 12232
rect 16482 12180 16488 12232
rect 16540 12180 16546 12232
rect 16577 12223 16635 12229
rect 16577 12189 16589 12223
rect 16623 12189 16635 12223
rect 16577 12183 16635 12189
rect 15286 12152 15292 12164
rect 14476 12124 15292 12152
rect 15286 12112 15292 12124
rect 15344 12112 15350 12164
rect 15930 12112 15936 12164
rect 15988 12152 15994 12164
rect 16592 12152 16620 12183
rect 16666 12180 16672 12232
rect 16724 12220 16730 12232
rect 16761 12223 16819 12229
rect 16761 12220 16773 12223
rect 16724 12192 16773 12220
rect 16724 12180 16730 12192
rect 16761 12189 16773 12192
rect 16807 12189 16819 12223
rect 16761 12183 16819 12189
rect 17034 12180 17040 12232
rect 17092 12180 17098 12232
rect 17512 12229 17540 12260
rect 17129 12223 17187 12229
rect 17129 12189 17141 12223
rect 17175 12189 17187 12223
rect 17129 12183 17187 12189
rect 17497 12223 17555 12229
rect 17497 12189 17509 12223
rect 17543 12189 17555 12223
rect 17497 12183 17555 12189
rect 17773 12223 17831 12229
rect 17773 12189 17785 12223
rect 17819 12189 17831 12223
rect 17773 12183 17831 12189
rect 18049 12223 18107 12229
rect 18049 12189 18061 12223
rect 18095 12189 18107 12223
rect 18049 12183 18107 12189
rect 15988 12124 16620 12152
rect 15988 12112 15994 12124
rect 14550 12084 14556 12096
rect 14108 12056 14556 12084
rect 14550 12044 14556 12056
rect 14608 12044 14614 12096
rect 14642 12044 14648 12096
rect 14700 12084 14706 12096
rect 17144 12084 17172 12183
rect 17788 12152 17816 12183
rect 18064 12152 18092 12183
rect 18138 12180 18144 12232
rect 18196 12180 18202 12232
rect 18524 12229 18552 12260
rect 18509 12223 18567 12229
rect 18509 12189 18521 12223
rect 18555 12220 18567 12223
rect 18966 12220 18972 12232
rect 18555 12192 18972 12220
rect 18555 12189 18567 12192
rect 18509 12183 18567 12189
rect 18966 12180 18972 12192
rect 19024 12180 19030 12232
rect 18598 12152 18604 12164
rect 17788 12124 18604 12152
rect 18598 12112 18604 12124
rect 18656 12112 18662 12164
rect 18138 12084 18144 12096
rect 14700 12056 18144 12084
rect 14700 12044 14706 12056
rect 18138 12044 18144 12056
rect 18196 12084 18202 12096
rect 19242 12084 19248 12096
rect 18196 12056 19248 12084
rect 18196 12044 18202 12056
rect 19242 12044 19248 12056
rect 19300 12044 19306 12096
rect 1104 11994 18860 12016
rect 1104 11942 2610 11994
rect 2662 11942 2674 11994
rect 2726 11942 2738 11994
rect 2790 11942 2802 11994
rect 2854 11942 2866 11994
rect 2918 11942 7610 11994
rect 7662 11942 7674 11994
rect 7726 11942 7738 11994
rect 7790 11942 7802 11994
rect 7854 11942 7866 11994
rect 7918 11942 12610 11994
rect 12662 11942 12674 11994
rect 12726 11942 12738 11994
rect 12790 11942 12802 11994
rect 12854 11942 12866 11994
rect 12918 11942 17610 11994
rect 17662 11942 17674 11994
rect 17726 11942 17738 11994
rect 17790 11942 17802 11994
rect 17854 11942 17866 11994
rect 17918 11942 18860 11994
rect 1104 11920 18860 11942
rect 1949 11883 2007 11889
rect 1949 11849 1961 11883
rect 1995 11880 2007 11883
rect 2498 11880 2504 11892
rect 1995 11852 2504 11880
rect 1995 11849 2007 11852
rect 1949 11843 2007 11849
rect 2498 11840 2504 11852
rect 2556 11840 2562 11892
rect 4062 11840 4068 11892
rect 4120 11880 4126 11892
rect 5258 11880 5264 11892
rect 4120 11852 5264 11880
rect 4120 11840 4126 11852
rect 5258 11840 5264 11852
rect 5316 11840 5322 11892
rect 5442 11840 5448 11892
rect 5500 11880 5506 11892
rect 5500 11852 6868 11880
rect 5500 11840 5506 11852
rect 1581 11815 1639 11821
rect 1581 11781 1593 11815
rect 1627 11781 1639 11815
rect 1581 11775 1639 11781
rect 1797 11815 1855 11821
rect 1797 11781 1809 11815
rect 1843 11812 1855 11815
rect 3418 11812 3424 11824
rect 1843 11784 3424 11812
rect 1843 11781 1855 11784
rect 1797 11775 1855 11781
rect 1596 11676 1624 11775
rect 3418 11772 3424 11784
rect 3476 11772 3482 11824
rect 3878 11772 3884 11824
rect 3936 11812 3942 11824
rect 5460 11812 5488 11840
rect 3936 11784 5488 11812
rect 3936 11772 3942 11784
rect 6362 11772 6368 11824
rect 6420 11812 6426 11824
rect 6840 11812 6868 11852
rect 7374 11840 7380 11892
rect 7432 11840 7438 11892
rect 7469 11883 7527 11889
rect 7469 11849 7481 11883
rect 7515 11880 7527 11883
rect 7558 11880 7564 11892
rect 7515 11852 7564 11880
rect 7515 11849 7527 11852
rect 7469 11843 7527 11849
rect 7558 11840 7564 11852
rect 7616 11880 7622 11892
rect 9766 11880 9772 11892
rect 7616 11852 9772 11880
rect 7616 11840 7622 11852
rect 9766 11840 9772 11852
rect 9824 11840 9830 11892
rect 10134 11880 10140 11892
rect 9968 11852 10140 11880
rect 7282 11812 7288 11824
rect 6420 11784 6776 11812
rect 6420 11772 6426 11784
rect 3050 11704 3056 11756
rect 3108 11704 3114 11756
rect 3602 11704 3608 11756
rect 3660 11744 3666 11756
rect 4154 11744 4160 11756
rect 3660 11716 4160 11744
rect 3660 11704 3666 11716
rect 4154 11704 4160 11716
rect 4212 11704 4218 11756
rect 4430 11704 4436 11756
rect 4488 11744 4494 11756
rect 4893 11747 4951 11753
rect 4893 11744 4905 11747
rect 4488 11716 4905 11744
rect 4488 11704 4494 11716
rect 4893 11713 4905 11716
rect 4939 11713 4951 11747
rect 4893 11707 4951 11713
rect 5166 11704 5172 11756
rect 5224 11704 5230 11756
rect 6748 11753 6776 11784
rect 6840 11784 7288 11812
rect 6840 11753 6868 11784
rect 7282 11772 7288 11784
rect 7340 11772 7346 11824
rect 9968 11812 9996 11852
rect 10134 11840 10140 11852
rect 10192 11840 10198 11892
rect 12802 11880 12808 11892
rect 10796 11852 12808 11880
rect 7484 11784 9996 11812
rect 6641 11747 6699 11753
rect 6641 11744 6653 11747
rect 5460 11716 6653 11744
rect 3510 11676 3516 11688
rect 1596 11648 3516 11676
rect 3510 11636 3516 11648
rect 3568 11676 3574 11688
rect 4246 11676 4252 11688
rect 3568 11648 4252 11676
rect 3568 11636 3574 11648
rect 4246 11636 4252 11648
rect 4304 11636 4310 11688
rect 2590 11568 2596 11620
rect 2648 11608 2654 11620
rect 4985 11611 5043 11617
rect 4985 11608 4997 11611
rect 2648 11580 4997 11608
rect 2648 11568 2654 11580
rect 4985 11577 4997 11580
rect 5031 11577 5043 11611
rect 4985 11571 5043 11577
rect 566 11500 572 11552
rect 624 11540 630 11552
rect 1486 11540 1492 11552
rect 624 11512 1492 11540
rect 624 11500 630 11512
rect 1486 11500 1492 11512
rect 1544 11500 1550 11552
rect 1765 11543 1823 11549
rect 1765 11509 1777 11543
rect 1811 11540 1823 11543
rect 1854 11540 1860 11552
rect 1811 11512 1860 11540
rect 1811 11509 1823 11512
rect 1765 11503 1823 11509
rect 1854 11500 1860 11512
rect 1912 11500 1918 11552
rect 2130 11500 2136 11552
rect 2188 11540 2194 11552
rect 2498 11540 2504 11552
rect 2188 11512 2504 11540
rect 2188 11500 2194 11512
rect 2498 11500 2504 11512
rect 2556 11500 2562 11552
rect 2866 11500 2872 11552
rect 2924 11540 2930 11552
rect 4706 11540 4712 11552
rect 2924 11512 4712 11540
rect 2924 11500 2930 11512
rect 4706 11500 4712 11512
rect 4764 11540 4770 11552
rect 5460 11540 5488 11716
rect 6641 11713 6653 11716
rect 6687 11713 6699 11747
rect 6641 11707 6699 11713
rect 6733 11747 6791 11753
rect 6733 11713 6745 11747
rect 6779 11713 6791 11747
rect 6733 11707 6791 11713
rect 6825 11747 6883 11753
rect 6825 11713 6837 11747
rect 6871 11713 6883 11747
rect 6825 11707 6883 11713
rect 7006 11704 7012 11756
rect 7064 11704 7070 11756
rect 7193 11747 7251 11753
rect 7193 11713 7205 11747
rect 7239 11744 7251 11747
rect 7374 11744 7380 11756
rect 7239 11716 7380 11744
rect 7239 11713 7251 11716
rect 7193 11707 7251 11713
rect 7374 11704 7380 11716
rect 7432 11704 7438 11756
rect 5629 11679 5687 11685
rect 5629 11645 5641 11679
rect 5675 11676 5687 11679
rect 7484 11676 7512 11784
rect 10042 11772 10048 11824
rect 10100 11812 10106 11824
rect 10796 11812 10824 11852
rect 12802 11840 12808 11852
rect 12860 11840 12866 11892
rect 13354 11840 13360 11892
rect 13412 11880 13418 11892
rect 13906 11880 13912 11892
rect 13412 11852 13912 11880
rect 13412 11840 13418 11852
rect 13906 11840 13912 11852
rect 13964 11840 13970 11892
rect 16482 11840 16488 11892
rect 16540 11880 16546 11892
rect 17034 11880 17040 11892
rect 16540 11852 17040 11880
rect 16540 11840 16546 11852
rect 17034 11840 17040 11852
rect 17092 11840 17098 11892
rect 10100 11784 10824 11812
rect 10100 11772 10106 11784
rect 10870 11772 10876 11824
rect 10928 11812 10934 11824
rect 10965 11815 11023 11821
rect 10965 11812 10977 11815
rect 10928 11784 10977 11812
rect 10928 11772 10934 11784
rect 10965 11781 10977 11784
rect 11011 11781 11023 11815
rect 10965 11775 11023 11781
rect 11054 11772 11060 11824
rect 11112 11812 11118 11824
rect 13722 11812 13728 11824
rect 11112 11784 13728 11812
rect 11112 11772 11118 11784
rect 13722 11772 13728 11784
rect 13780 11772 13786 11824
rect 15470 11772 15476 11824
rect 15528 11812 15534 11824
rect 16574 11812 16580 11824
rect 15528 11784 16580 11812
rect 15528 11772 15534 11784
rect 16574 11772 16580 11784
rect 16632 11772 16638 11824
rect 16850 11772 16856 11824
rect 16908 11812 16914 11824
rect 16908 11784 17816 11812
rect 16908 11772 16914 11784
rect 7561 11747 7619 11753
rect 7561 11713 7573 11747
rect 7607 11713 7619 11747
rect 7561 11707 7619 11713
rect 5675 11648 7512 11676
rect 5675 11645 5687 11648
rect 5629 11639 5687 11645
rect 6086 11568 6092 11620
rect 6144 11608 6150 11620
rect 6454 11608 6460 11620
rect 6144 11580 6460 11608
rect 6144 11568 6150 11580
rect 6454 11568 6460 11580
rect 6512 11568 6518 11620
rect 6546 11568 6552 11620
rect 6604 11608 6610 11620
rect 6730 11608 6736 11620
rect 6604 11580 6736 11608
rect 6604 11568 6610 11580
rect 6730 11568 6736 11580
rect 6788 11608 6794 11620
rect 7576 11608 7604 11707
rect 7742 11704 7748 11756
rect 7800 11744 7806 11756
rect 8386 11744 8392 11756
rect 7800 11716 8392 11744
rect 7800 11704 7806 11716
rect 8386 11704 8392 11716
rect 8444 11704 8450 11756
rect 9490 11704 9496 11756
rect 9548 11744 9554 11756
rect 9585 11747 9643 11753
rect 9585 11744 9597 11747
rect 9548 11716 9597 11744
rect 9548 11704 9554 11716
rect 9585 11713 9597 11716
rect 9631 11713 9643 11747
rect 9585 11707 9643 11713
rect 9674 11704 9680 11756
rect 9732 11744 9738 11756
rect 9769 11747 9827 11753
rect 9769 11744 9781 11747
rect 9732 11716 9781 11744
rect 9732 11704 9738 11716
rect 9769 11713 9781 11716
rect 9815 11744 9827 11747
rect 9815 11716 10456 11744
rect 9815 11713 9827 11716
rect 9769 11707 9827 11713
rect 7834 11636 7840 11688
rect 7892 11636 7898 11688
rect 8018 11636 8024 11688
rect 8076 11636 8082 11688
rect 8113 11679 8171 11685
rect 8113 11645 8125 11679
rect 8159 11676 8171 11679
rect 8481 11679 8539 11685
rect 8159 11648 8432 11676
rect 8159 11645 8171 11648
rect 8113 11639 8171 11645
rect 7852 11608 7880 11636
rect 8404 11620 8432 11648
rect 8481 11645 8493 11679
rect 8527 11645 8539 11679
rect 8481 11639 8539 11645
rect 6788 11580 7604 11608
rect 7656 11580 7880 11608
rect 6788 11568 6794 11580
rect 4764 11512 5488 11540
rect 4764 11500 4770 11512
rect 5534 11500 5540 11552
rect 5592 11540 5598 11552
rect 5718 11540 5724 11552
rect 5592 11512 5724 11540
rect 5592 11500 5598 11512
rect 5718 11500 5724 11512
rect 5776 11500 5782 11552
rect 6362 11500 6368 11552
rect 6420 11500 6426 11552
rect 6472 11540 6500 11568
rect 7656 11540 7684 11580
rect 8386 11568 8392 11620
rect 8444 11568 8450 11620
rect 8496 11608 8524 11639
rect 9950 11636 9956 11688
rect 10008 11676 10014 11688
rect 10428 11676 10456 11716
rect 10502 11704 10508 11756
rect 10560 11744 10566 11756
rect 10778 11744 10784 11756
rect 10560 11716 10784 11744
rect 10560 11704 10566 11716
rect 10778 11704 10784 11716
rect 10836 11704 10842 11756
rect 11146 11704 11152 11756
rect 11204 11704 11210 11756
rect 11256 11753 11468 11754
rect 11241 11747 11468 11753
rect 11241 11713 11253 11747
rect 11287 11744 11468 11747
rect 11514 11744 11520 11756
rect 11287 11726 11520 11744
rect 11287 11713 11299 11726
rect 11440 11716 11520 11726
rect 11241 11707 11299 11713
rect 11514 11704 11520 11716
rect 11572 11704 11578 11756
rect 12802 11704 12808 11756
rect 12860 11744 12866 11756
rect 13909 11747 13967 11753
rect 13909 11744 13921 11747
rect 12860 11716 13921 11744
rect 12860 11704 12866 11716
rect 13909 11713 13921 11716
rect 13955 11713 13967 11747
rect 14553 11747 14611 11753
rect 14553 11744 14565 11747
rect 13909 11707 13967 11713
rect 14016 11716 14565 11744
rect 14016 11688 14044 11716
rect 14553 11713 14565 11716
rect 14599 11713 14611 11747
rect 14553 11707 14611 11713
rect 17402 11704 17408 11756
rect 17460 11704 17466 11756
rect 17788 11753 17816 11784
rect 18230 11772 18236 11824
rect 18288 11772 18294 11824
rect 17589 11747 17647 11753
rect 17589 11713 17601 11747
rect 17635 11713 17647 11747
rect 17589 11707 17647 11713
rect 17773 11747 17831 11753
rect 17773 11713 17785 11747
rect 17819 11713 17831 11747
rect 17773 11707 17831 11713
rect 10008 11648 10180 11676
rect 10428 11648 11928 11676
rect 10008 11636 10014 11648
rect 8938 11608 8944 11620
rect 8496 11580 8944 11608
rect 8938 11568 8944 11580
rect 8996 11568 9002 11620
rect 9677 11611 9735 11617
rect 9677 11577 9689 11611
rect 9723 11608 9735 11611
rect 10042 11608 10048 11620
rect 9723 11580 10048 11608
rect 9723 11577 9735 11580
rect 9677 11571 9735 11577
rect 10042 11568 10048 11580
rect 10100 11568 10106 11620
rect 10152 11608 10180 11648
rect 11057 11611 11115 11617
rect 11057 11608 11069 11611
rect 10152 11580 11069 11608
rect 11057 11577 11069 11580
rect 11103 11577 11115 11611
rect 11057 11571 11115 11577
rect 11422 11568 11428 11620
rect 11480 11608 11486 11620
rect 11790 11608 11796 11620
rect 11480 11580 11796 11608
rect 11480 11568 11486 11580
rect 11790 11568 11796 11580
rect 11848 11568 11854 11620
rect 11900 11608 11928 11648
rect 12342 11636 12348 11688
rect 12400 11676 12406 11688
rect 13817 11679 13875 11685
rect 13817 11676 13829 11679
rect 12400 11648 13829 11676
rect 12400 11636 12406 11648
rect 13817 11645 13829 11648
rect 13863 11645 13875 11679
rect 13817 11639 13875 11645
rect 13998 11636 14004 11688
rect 14056 11636 14062 11688
rect 14366 11636 14372 11688
rect 14424 11636 14430 11688
rect 14461 11679 14519 11685
rect 14461 11645 14473 11679
rect 14507 11645 14519 11679
rect 14461 11639 14519 11645
rect 13262 11608 13268 11620
rect 11900 11580 13268 11608
rect 13262 11568 13268 11580
rect 13320 11568 13326 11620
rect 14476 11608 14504 11639
rect 14642 11636 14648 11688
rect 14700 11636 14706 11688
rect 15930 11636 15936 11688
rect 15988 11676 15994 11688
rect 16758 11676 16764 11688
rect 15988 11648 16764 11676
rect 15988 11636 15994 11648
rect 16758 11636 16764 11648
rect 16816 11636 16822 11688
rect 17604 11676 17632 11707
rect 18506 11676 18512 11688
rect 17604 11648 18512 11676
rect 18506 11636 18512 11648
rect 18564 11636 18570 11688
rect 14826 11608 14832 11620
rect 14476 11580 14832 11608
rect 14826 11568 14832 11580
rect 14884 11568 14890 11620
rect 6472 11512 7684 11540
rect 7837 11543 7895 11549
rect 7837 11509 7849 11543
rect 7883 11540 7895 11543
rect 7926 11540 7932 11552
rect 7883 11512 7932 11540
rect 7883 11509 7895 11512
rect 7837 11503 7895 11509
rect 7926 11500 7932 11512
rect 7984 11500 7990 11552
rect 8570 11500 8576 11552
rect 8628 11540 8634 11552
rect 13541 11543 13599 11549
rect 13541 11540 13553 11543
rect 8628 11512 13553 11540
rect 8628 11500 8634 11512
rect 13541 11509 13553 11512
rect 13587 11509 13599 11543
rect 13541 11503 13599 11509
rect 13722 11500 13728 11552
rect 13780 11540 13786 11552
rect 14185 11543 14243 11549
rect 14185 11540 14197 11543
rect 13780 11512 14197 11540
rect 13780 11500 13786 11512
rect 14185 11509 14197 11512
rect 14231 11509 14243 11543
rect 14185 11503 14243 11509
rect 15838 11500 15844 11552
rect 15896 11540 15902 11552
rect 16758 11540 16764 11552
rect 15896 11512 16764 11540
rect 15896 11500 15902 11512
rect 16758 11500 16764 11512
rect 16816 11540 16822 11552
rect 17494 11540 17500 11552
rect 16816 11512 17500 11540
rect 16816 11500 16822 11512
rect 17494 11500 17500 11512
rect 17552 11500 17558 11552
rect 1104 11450 18860 11472
rect 1104 11398 1950 11450
rect 2002 11398 2014 11450
rect 2066 11398 2078 11450
rect 2130 11398 2142 11450
rect 2194 11398 2206 11450
rect 2258 11398 6950 11450
rect 7002 11398 7014 11450
rect 7066 11398 7078 11450
rect 7130 11398 7142 11450
rect 7194 11398 7206 11450
rect 7258 11398 11950 11450
rect 12002 11398 12014 11450
rect 12066 11398 12078 11450
rect 12130 11398 12142 11450
rect 12194 11398 12206 11450
rect 12258 11398 16950 11450
rect 17002 11398 17014 11450
rect 17066 11398 17078 11450
rect 17130 11398 17142 11450
rect 17194 11398 17206 11450
rect 17258 11398 18860 11450
rect 1104 11376 18860 11398
rect 1394 11296 1400 11348
rect 1452 11296 1458 11348
rect 2222 11296 2228 11348
rect 2280 11336 2286 11348
rect 2590 11336 2596 11348
rect 2280 11308 2596 11336
rect 2280 11296 2286 11308
rect 2590 11296 2596 11308
rect 2648 11296 2654 11348
rect 3694 11296 3700 11348
rect 3752 11336 3758 11348
rect 4154 11336 4160 11348
rect 3752 11308 4160 11336
rect 3752 11296 3758 11308
rect 4154 11296 4160 11308
rect 4212 11296 4218 11348
rect 4614 11296 4620 11348
rect 4672 11336 4678 11348
rect 4709 11339 4767 11345
rect 4709 11336 4721 11339
rect 4672 11308 4721 11336
rect 4672 11296 4678 11308
rect 4709 11305 4721 11308
rect 4755 11305 4767 11339
rect 5537 11339 5595 11345
rect 5537 11336 5549 11339
rect 4709 11299 4767 11305
rect 4816 11308 5549 11336
rect 1412 11200 1440 11296
rect 1578 11228 1584 11280
rect 1636 11268 1642 11280
rect 2958 11268 2964 11280
rect 1636 11240 2964 11268
rect 1636 11228 1642 11240
rect 2958 11228 2964 11240
rect 3016 11228 3022 11280
rect 4062 11228 4068 11280
rect 4120 11268 4126 11280
rect 4430 11268 4436 11280
rect 4120 11240 4436 11268
rect 4120 11228 4126 11240
rect 4430 11228 4436 11240
rect 4488 11228 4494 11280
rect 1320 11172 1440 11200
rect 1320 11064 1348 11172
rect 1486 11160 1492 11212
rect 1544 11200 1550 11212
rect 1762 11200 1768 11212
rect 1544 11172 1768 11200
rect 1544 11160 1550 11172
rect 1762 11160 1768 11172
rect 1820 11160 1826 11212
rect 4614 11160 4620 11212
rect 4672 11200 4678 11212
rect 4816 11200 4844 11308
rect 5537 11305 5549 11308
rect 5583 11305 5595 11339
rect 5537 11299 5595 11305
rect 5994 11296 6000 11348
rect 6052 11336 6058 11348
rect 6089 11339 6147 11345
rect 6089 11336 6101 11339
rect 6052 11308 6101 11336
rect 6052 11296 6058 11308
rect 6089 11305 6101 11308
rect 6135 11305 6147 11339
rect 6089 11299 6147 11305
rect 6730 11296 6736 11348
rect 6788 11336 6794 11348
rect 7098 11336 7104 11348
rect 6788 11308 7104 11336
rect 6788 11296 6794 11308
rect 7098 11296 7104 11308
rect 7156 11296 7162 11348
rect 10870 11336 10876 11348
rect 7579 11308 9628 11336
rect 7579 11268 7607 11308
rect 4672 11172 4844 11200
rect 4908 11240 7607 11268
rect 7653 11271 7711 11277
rect 4672 11160 4678 11172
rect 1394 11092 1400 11144
rect 1452 11092 1458 11144
rect 3878 11092 3884 11144
rect 3936 11132 3942 11144
rect 3973 11135 4031 11141
rect 3973 11132 3985 11135
rect 3936 11104 3985 11132
rect 3936 11092 3942 11104
rect 3973 11101 3985 11104
rect 4019 11101 4031 11135
rect 3973 11095 4031 11101
rect 4525 11135 4583 11141
rect 4525 11101 4537 11135
rect 4571 11132 4583 11135
rect 4908 11132 4936 11240
rect 7653 11237 7665 11271
rect 7699 11268 7711 11271
rect 8110 11268 8116 11280
rect 7699 11240 8116 11268
rect 7699 11237 7711 11240
rect 7653 11231 7711 11237
rect 8110 11228 8116 11240
rect 8168 11228 8174 11280
rect 9600 11268 9628 11308
rect 9968 11308 10876 11336
rect 9968 11268 9996 11308
rect 10870 11296 10876 11308
rect 10928 11336 10934 11348
rect 14182 11336 14188 11348
rect 10928 11308 14188 11336
rect 10928 11296 10934 11308
rect 14182 11296 14188 11308
rect 14240 11296 14246 11348
rect 14734 11296 14740 11348
rect 14792 11336 14798 11348
rect 16942 11336 16948 11348
rect 14792 11308 16948 11336
rect 14792 11296 14798 11308
rect 16942 11296 16948 11308
rect 17000 11296 17006 11348
rect 9600 11240 9996 11268
rect 10778 11228 10784 11280
rect 10836 11268 10842 11280
rect 10836 11240 12664 11268
rect 10836 11228 10842 11240
rect 5261 11203 5319 11209
rect 5261 11169 5273 11203
rect 5307 11200 5319 11203
rect 5718 11200 5724 11212
rect 5307 11172 5724 11200
rect 5307 11169 5319 11172
rect 5261 11163 5319 11169
rect 5718 11160 5724 11172
rect 5776 11200 5782 11212
rect 6914 11200 6920 11212
rect 5776 11172 6132 11200
rect 5776 11160 5782 11172
rect 4571 11104 4936 11132
rect 4571 11101 4583 11104
rect 4525 11095 4583 11101
rect 5074 11092 5080 11144
rect 5132 11092 5138 11144
rect 5442 11142 5448 11144
rect 5368 11141 5448 11142
rect 5353 11135 5448 11141
rect 5353 11132 5365 11135
rect 5184 11104 5365 11132
rect 1673 11067 1731 11073
rect 1320 11036 1440 11064
rect 1412 11008 1440 11036
rect 1673 11033 1685 11067
rect 1719 11064 1731 11067
rect 1762 11064 1768 11076
rect 1719 11036 1768 11064
rect 1719 11033 1731 11036
rect 1673 11027 1731 11033
rect 1762 11024 1768 11036
rect 1820 11064 1826 11076
rect 3050 11064 3056 11076
rect 1820 11036 3056 11064
rect 1820 11024 1826 11036
rect 3050 11024 3056 11036
rect 3108 11064 3114 11076
rect 4798 11064 4804 11076
rect 3108 11036 4804 11064
rect 3108 11024 3114 11036
rect 4798 11024 4804 11036
rect 4856 11064 4862 11076
rect 5184 11064 5212 11104
rect 5353 11101 5365 11104
rect 5399 11114 5448 11135
rect 5399 11101 5411 11114
rect 5353 11095 5411 11101
rect 5442 11092 5448 11114
rect 5500 11092 5506 11144
rect 5994 11092 6000 11144
rect 6052 11092 6058 11144
rect 4856 11036 5212 11064
rect 6104 11064 6132 11172
rect 6288 11172 6920 11200
rect 6178 11092 6184 11144
rect 6236 11141 6242 11144
rect 6236 11132 6247 11141
rect 6288 11132 6316 11172
rect 6914 11160 6920 11172
rect 6972 11160 6978 11212
rect 7098 11160 7104 11212
rect 7156 11200 7162 11212
rect 7285 11203 7343 11209
rect 7285 11200 7297 11203
rect 7156 11172 7297 11200
rect 7156 11160 7162 11172
rect 7285 11169 7297 11172
rect 7331 11169 7343 11203
rect 7285 11163 7343 11169
rect 7466 11160 7472 11212
rect 7524 11200 7530 11212
rect 7745 11203 7803 11209
rect 7745 11200 7757 11203
rect 7524 11172 7757 11200
rect 7524 11160 7530 11172
rect 7745 11169 7757 11172
rect 7791 11169 7803 11203
rect 7745 11163 7803 11169
rect 8570 11160 8576 11212
rect 8628 11200 8634 11212
rect 8754 11200 8760 11212
rect 8628 11172 8760 11200
rect 8628 11160 8634 11172
rect 8754 11160 8760 11172
rect 8812 11160 8818 11212
rect 9490 11160 9496 11212
rect 9548 11200 9554 11212
rect 10137 11203 10195 11209
rect 9548 11172 10088 11200
rect 9548 11160 9554 11172
rect 10060 11144 10088 11172
rect 10137 11169 10149 11203
rect 10183 11200 10195 11203
rect 10318 11200 10324 11212
rect 10183 11172 10324 11200
rect 10183 11169 10195 11172
rect 10137 11163 10195 11169
rect 10318 11160 10324 11172
rect 10376 11200 10382 11212
rect 10597 11203 10655 11209
rect 10597 11200 10609 11203
rect 10376 11172 10609 11200
rect 10376 11160 10382 11172
rect 10597 11169 10609 11172
rect 10643 11169 10655 11203
rect 10597 11163 10655 11169
rect 10704 11172 11100 11200
rect 6236 11104 6316 11132
rect 6236 11095 6247 11104
rect 6236 11092 6242 11095
rect 6822 11092 6828 11144
rect 6880 11132 6886 11144
rect 6880 11104 9812 11132
rect 6880 11092 6886 11104
rect 6104 11036 6868 11064
rect 4856 11024 4862 11036
rect 1394 10956 1400 11008
rect 1452 10956 1458 11008
rect 3418 10956 3424 11008
rect 3476 10996 3482 11008
rect 6730 10996 6736 11008
rect 3476 10968 6736 10996
rect 3476 10956 3482 10968
rect 6730 10956 6736 10968
rect 6788 10956 6794 11008
rect 6840 10996 6868 11036
rect 7006 11024 7012 11076
rect 7064 11064 7070 11076
rect 7742 11064 7748 11076
rect 7064 11036 7748 11064
rect 7064 11024 7070 11036
rect 7742 11024 7748 11036
rect 7800 11024 7806 11076
rect 7834 11024 7840 11076
rect 7892 11064 7898 11076
rect 8938 11064 8944 11076
rect 7892 11036 8944 11064
rect 7892 11024 7898 11036
rect 8938 11024 8944 11036
rect 8996 11024 9002 11076
rect 9214 11024 9220 11076
rect 9272 11024 9278 11076
rect 9784 11064 9812 11104
rect 10042 11092 10048 11144
rect 10100 11092 10106 11144
rect 10704 11064 10732 11172
rect 10781 11135 10839 11141
rect 10781 11101 10793 11135
rect 10827 11101 10839 11135
rect 10781 11095 10839 11101
rect 9784 11036 10732 11064
rect 10796 11064 10824 11095
rect 10962 11092 10968 11144
rect 11020 11092 11026 11144
rect 11072 11141 11100 11172
rect 11238 11160 11244 11212
rect 11296 11200 11302 11212
rect 12526 11200 12532 11212
rect 11296 11172 12532 11200
rect 11296 11160 11302 11172
rect 12526 11160 12532 11172
rect 12584 11160 12590 11212
rect 12636 11200 12664 11240
rect 12710 11228 12716 11280
rect 12768 11268 12774 11280
rect 13814 11268 13820 11280
rect 12768 11240 13820 11268
rect 12768 11228 12774 11240
rect 13814 11228 13820 11240
rect 13872 11228 13878 11280
rect 15838 11228 15844 11280
rect 15896 11228 15902 11280
rect 16393 11271 16451 11277
rect 16393 11237 16405 11271
rect 16439 11268 16451 11271
rect 17954 11268 17960 11280
rect 16439 11240 17960 11268
rect 16439 11237 16451 11240
rect 16393 11231 16451 11237
rect 17954 11228 17960 11240
rect 18012 11228 18018 11280
rect 12636 11172 16712 11200
rect 11057 11135 11115 11141
rect 11057 11101 11069 11135
rect 11103 11132 11115 11135
rect 11698 11132 11704 11144
rect 11103 11104 11704 11132
rect 11103 11101 11115 11104
rect 11057 11095 11115 11101
rect 11698 11092 11704 11104
rect 11756 11132 11762 11144
rect 11756 11104 11836 11132
rect 11756 11092 11762 11104
rect 11808 11064 11836 11104
rect 11882 11092 11888 11144
rect 11940 11132 11946 11144
rect 12710 11132 12716 11144
rect 11940 11104 12716 11132
rect 11940 11092 11946 11104
rect 12710 11092 12716 11104
rect 12768 11092 12774 11144
rect 13170 11092 13176 11144
rect 13228 11092 13234 11144
rect 14366 11092 14372 11144
rect 14424 11132 14430 11144
rect 15654 11132 15660 11144
rect 14424 11104 15660 11132
rect 14424 11092 14430 11104
rect 15654 11092 15660 11104
rect 15712 11092 15718 11144
rect 15838 11092 15844 11144
rect 15896 11132 15902 11144
rect 16684 11141 16712 11172
rect 16850 11160 16856 11212
rect 16908 11160 16914 11212
rect 16209 11135 16267 11141
rect 16209 11132 16221 11135
rect 15896 11104 16221 11132
rect 15896 11092 15902 11104
rect 16209 11101 16221 11104
rect 16255 11101 16267 11135
rect 16209 11095 16267 11101
rect 16669 11135 16727 11141
rect 16669 11101 16681 11135
rect 16715 11101 16727 11135
rect 16669 11095 16727 11101
rect 17037 11135 17095 11141
rect 17037 11101 17049 11135
rect 17083 11101 17095 11135
rect 17037 11095 17095 11101
rect 11974 11064 11980 11076
rect 10796 11036 11744 11064
rect 11808 11036 11980 11064
rect 9490 10996 9496 11008
rect 6840 10968 9496 10996
rect 9490 10956 9496 10968
rect 9548 10956 9554 11008
rect 10042 10956 10048 11008
rect 10100 10996 10106 11008
rect 11606 10996 11612 11008
rect 10100 10968 11612 10996
rect 10100 10956 10106 10968
rect 11606 10956 11612 10968
rect 11664 10956 11670 11008
rect 11716 10996 11744 11036
rect 11974 11024 11980 11036
rect 12032 11024 12038 11076
rect 12434 11024 12440 11076
rect 12492 11064 12498 11076
rect 13188 11064 13216 11092
rect 12492 11036 13216 11064
rect 12492 11024 12498 11036
rect 16482 11024 16488 11076
rect 16540 11064 16546 11076
rect 17052 11064 17080 11095
rect 17494 11092 17500 11144
rect 17552 11092 17558 11144
rect 17770 11092 17776 11144
rect 17828 11092 17834 11144
rect 18046 11092 18052 11144
rect 18104 11132 18110 11144
rect 18141 11135 18199 11141
rect 18141 11132 18153 11135
rect 18104 11104 18153 11132
rect 18104 11092 18110 11104
rect 18141 11101 18153 11104
rect 18187 11101 18199 11135
rect 18141 11095 18199 11101
rect 16540 11036 17080 11064
rect 16540 11024 16546 11036
rect 17402 11024 17408 11076
rect 17460 11064 17466 11076
rect 18064 11064 18092 11092
rect 17460 11036 18092 11064
rect 17460 11024 17466 11036
rect 12158 10996 12164 11008
rect 11716 10968 12164 10996
rect 12158 10956 12164 10968
rect 12216 10956 12222 11008
rect 15102 10956 15108 11008
rect 15160 10996 15166 11008
rect 15562 10996 15568 11008
rect 15160 10968 15568 10996
rect 15160 10956 15166 10968
rect 15562 10956 15568 10968
rect 15620 10956 15626 11008
rect 17862 10956 17868 11008
rect 17920 10996 17926 11008
rect 18690 10996 18696 11008
rect 17920 10968 18696 10996
rect 17920 10956 17926 10968
rect 18690 10956 18696 10968
rect 18748 10956 18754 11008
rect 1104 10906 18860 10928
rect 1104 10854 2610 10906
rect 2662 10854 2674 10906
rect 2726 10854 2738 10906
rect 2790 10854 2802 10906
rect 2854 10854 2866 10906
rect 2918 10854 7610 10906
rect 7662 10854 7674 10906
rect 7726 10854 7738 10906
rect 7790 10854 7802 10906
rect 7854 10854 7866 10906
rect 7918 10854 12610 10906
rect 12662 10854 12674 10906
rect 12726 10854 12738 10906
rect 12790 10854 12802 10906
rect 12854 10854 12866 10906
rect 12918 10854 17610 10906
rect 17662 10854 17674 10906
rect 17726 10854 17738 10906
rect 17790 10854 17802 10906
rect 17854 10854 17866 10906
rect 17918 10854 18860 10906
rect 1104 10832 18860 10854
rect 2222 10752 2228 10804
rect 2280 10792 2286 10804
rect 2590 10792 2596 10804
rect 2280 10764 2596 10792
rect 2280 10752 2286 10764
rect 2590 10752 2596 10764
rect 2648 10752 2654 10804
rect 3418 10752 3424 10804
rect 3476 10792 3482 10804
rect 3602 10792 3608 10804
rect 3476 10764 3608 10792
rect 3476 10752 3482 10764
rect 3602 10752 3608 10764
rect 3660 10752 3666 10804
rect 4338 10752 4344 10804
rect 4396 10792 4402 10804
rect 4433 10795 4491 10801
rect 4433 10792 4445 10795
rect 4396 10764 4445 10792
rect 4396 10752 4402 10764
rect 4433 10761 4445 10764
rect 4479 10792 4491 10795
rect 4890 10792 4896 10804
rect 4479 10764 4896 10792
rect 4479 10761 4491 10764
rect 4433 10755 4491 10761
rect 4890 10752 4896 10764
rect 4948 10752 4954 10804
rect 4982 10752 4988 10804
rect 5040 10752 5046 10804
rect 5350 10752 5356 10804
rect 5408 10752 5414 10804
rect 5442 10752 5448 10804
rect 5500 10792 5506 10804
rect 8202 10792 8208 10804
rect 5500 10764 8208 10792
rect 5500 10752 5506 10764
rect 8202 10752 8208 10764
rect 8260 10752 8266 10804
rect 11790 10792 11796 10804
rect 8772 10764 11796 10792
rect 2866 10684 2872 10736
rect 2924 10724 2930 10736
rect 4706 10724 4712 10736
rect 2924 10696 4712 10724
rect 2924 10684 2930 10696
rect 4706 10684 4712 10696
rect 4764 10684 4770 10736
rect 4798 10684 4804 10736
rect 4856 10724 4862 10736
rect 5000 10724 5028 10752
rect 5368 10724 5396 10752
rect 7834 10724 7840 10736
rect 4856 10696 5028 10724
rect 5184 10696 5948 10724
rect 4856 10684 4862 10696
rect 3053 10659 3111 10665
rect 3053 10625 3065 10659
rect 3099 10656 3111 10659
rect 3602 10656 3608 10668
rect 3099 10628 3608 10656
rect 3099 10625 3111 10628
rect 3053 10619 3111 10625
rect 3602 10616 3608 10628
rect 3660 10616 3666 10668
rect 3970 10616 3976 10668
rect 4028 10616 4034 10668
rect 4338 10616 4344 10668
rect 4396 10656 4402 10668
rect 4436 10659 4494 10665
rect 4436 10656 4448 10659
rect 4396 10628 4448 10656
rect 4396 10616 4402 10628
rect 4436 10625 4448 10628
rect 4482 10625 4494 10659
rect 4436 10619 4494 10625
rect 5184 10600 5212 10696
rect 5721 10659 5779 10665
rect 5721 10625 5733 10659
rect 5767 10625 5779 10659
rect 5721 10619 5779 10625
rect 5813 10659 5871 10665
rect 5813 10625 5825 10659
rect 5859 10654 5871 10659
rect 5920 10654 5948 10696
rect 6932 10696 7840 10724
rect 5859 10626 5948 10654
rect 5859 10625 5871 10626
rect 5813 10619 5871 10625
rect 3329 10591 3387 10597
rect 3329 10557 3341 10591
rect 3375 10588 3387 10591
rect 4246 10588 4252 10600
rect 3375 10560 4252 10588
rect 3375 10557 3387 10560
rect 3329 10551 3387 10557
rect 4246 10548 4252 10560
rect 4304 10548 4310 10600
rect 5166 10548 5172 10600
rect 5224 10548 5230 10600
rect 5258 10548 5264 10600
rect 5316 10588 5322 10600
rect 5353 10591 5411 10597
rect 5353 10588 5365 10591
rect 5316 10560 5365 10588
rect 5316 10548 5322 10560
rect 5353 10557 5365 10560
rect 5399 10557 5411 10591
rect 5353 10551 5411 10557
rect 5442 10548 5448 10600
rect 5500 10548 5506 10600
rect 5736 10588 5764 10619
rect 5994 10616 6000 10668
rect 6052 10656 6058 10668
rect 6052 10628 6232 10656
rect 6052 10616 6058 10628
rect 6086 10588 6092 10600
rect 5736 10560 6092 10588
rect 6086 10548 6092 10560
rect 6144 10548 6150 10600
rect 6204 10588 6232 10628
rect 6270 10616 6276 10668
rect 6328 10656 6334 10668
rect 6365 10659 6423 10665
rect 6365 10656 6377 10659
rect 6328 10628 6377 10656
rect 6328 10616 6334 10628
rect 6365 10625 6377 10628
rect 6411 10625 6423 10659
rect 6365 10619 6423 10625
rect 6733 10659 6791 10665
rect 6733 10625 6745 10659
rect 6779 10656 6791 10659
rect 6822 10656 6828 10668
rect 6779 10628 6828 10656
rect 6779 10625 6791 10628
rect 6733 10619 6791 10625
rect 6822 10616 6828 10628
rect 6880 10616 6886 10668
rect 6932 10665 6960 10696
rect 7834 10684 7840 10696
rect 7892 10684 7898 10736
rect 8772 10724 8800 10764
rect 11790 10752 11796 10764
rect 11848 10752 11854 10804
rect 12618 10752 12624 10804
rect 12676 10792 12682 10804
rect 13262 10792 13268 10804
rect 12676 10764 13268 10792
rect 12676 10752 12682 10764
rect 13262 10752 13268 10764
rect 13320 10752 13326 10804
rect 13630 10752 13636 10804
rect 13688 10792 13694 10804
rect 13725 10795 13783 10801
rect 13725 10792 13737 10795
rect 13688 10764 13737 10792
rect 13688 10752 13694 10764
rect 13725 10761 13737 10764
rect 13771 10761 13783 10795
rect 13725 10755 13783 10761
rect 14182 10752 14188 10804
rect 14240 10792 14246 10804
rect 14240 10764 14412 10792
rect 14240 10752 14246 10764
rect 7944 10696 8800 10724
rect 6917 10659 6975 10665
rect 6917 10625 6929 10659
rect 6963 10625 6975 10659
rect 6917 10619 6975 10625
rect 7190 10616 7196 10668
rect 7248 10616 7254 10668
rect 7282 10616 7288 10668
rect 7340 10616 7346 10668
rect 7650 10616 7656 10668
rect 7708 10656 7714 10668
rect 7944 10656 7972 10696
rect 9490 10684 9496 10736
rect 9548 10724 9554 10736
rect 9766 10724 9772 10736
rect 9548 10696 9772 10724
rect 9548 10684 9554 10696
rect 9766 10684 9772 10696
rect 9824 10684 9830 10736
rect 9950 10684 9956 10736
rect 10008 10724 10014 10736
rect 11882 10724 11888 10736
rect 10008 10696 11888 10724
rect 10008 10684 10014 10696
rect 11882 10684 11888 10696
rect 11940 10684 11946 10736
rect 11992 10696 14320 10724
rect 7708 10628 7972 10656
rect 7708 10616 7714 10628
rect 8202 10616 8208 10668
rect 8260 10656 8266 10668
rect 11054 10656 11060 10668
rect 8260 10628 11060 10656
rect 8260 10616 8266 10628
rect 11054 10616 11060 10628
rect 11112 10616 11118 10668
rect 11514 10656 11520 10668
rect 11164 10628 11520 10656
rect 7466 10588 7472 10600
rect 6204 10560 7472 10588
rect 7466 10548 7472 10560
rect 7524 10548 7530 10600
rect 7742 10548 7748 10600
rect 7800 10588 7806 10600
rect 11164 10588 11192 10628
rect 11514 10616 11520 10628
rect 11572 10616 11578 10668
rect 11606 10616 11612 10668
rect 11664 10616 11670 10668
rect 11790 10616 11796 10668
rect 11848 10616 11854 10668
rect 11992 10588 12020 10696
rect 12158 10616 12164 10668
rect 12216 10656 12222 10668
rect 12710 10656 12716 10668
rect 12216 10628 12716 10656
rect 12216 10616 12222 10628
rect 12710 10616 12716 10628
rect 12768 10616 12774 10668
rect 12894 10616 12900 10668
rect 12952 10656 12958 10668
rect 13265 10659 13323 10665
rect 13265 10656 13277 10659
rect 12952 10628 13277 10656
rect 12952 10616 12958 10628
rect 13265 10625 13277 10628
rect 13311 10625 13323 10659
rect 13265 10619 13323 10625
rect 13449 10659 13507 10665
rect 13449 10625 13461 10659
rect 13495 10656 13507 10659
rect 13909 10659 13967 10665
rect 13495 10628 13584 10656
rect 13495 10625 13507 10628
rect 13449 10619 13507 10625
rect 13556 10600 13584 10628
rect 13909 10625 13921 10659
rect 13955 10625 13967 10659
rect 13909 10619 13967 10625
rect 7800 10560 11192 10588
rect 11256 10560 12020 10588
rect 7800 10548 7806 10560
rect 3605 10523 3663 10529
rect 3605 10489 3617 10523
rect 3651 10520 3663 10523
rect 3970 10520 3976 10532
rect 3651 10492 3976 10520
rect 3651 10489 3663 10492
rect 3605 10483 3663 10489
rect 3970 10480 3976 10492
rect 4028 10480 4034 10532
rect 4617 10523 4675 10529
rect 4617 10489 4629 10523
rect 4663 10520 4675 10523
rect 5902 10520 5908 10532
rect 4663 10492 5908 10520
rect 4663 10489 4675 10492
rect 4617 10483 4675 10489
rect 5902 10480 5908 10492
rect 5960 10480 5966 10532
rect 5994 10480 6000 10532
rect 6052 10480 6058 10532
rect 6641 10523 6699 10529
rect 6641 10520 6653 10523
rect 6104 10492 6653 10520
rect 3421 10455 3479 10461
rect 3421 10421 3433 10455
rect 3467 10452 3479 10455
rect 3510 10452 3516 10464
rect 3467 10424 3516 10452
rect 3467 10421 3479 10424
rect 3421 10415 3479 10421
rect 3510 10412 3516 10424
rect 3568 10412 3574 10464
rect 3694 10412 3700 10464
rect 3752 10452 3758 10464
rect 4065 10455 4123 10461
rect 4065 10452 4077 10455
rect 3752 10424 4077 10452
rect 3752 10412 3758 10424
rect 4065 10421 4077 10424
rect 4111 10421 4123 10455
rect 4065 10415 4123 10421
rect 5718 10412 5724 10464
rect 5776 10452 5782 10464
rect 6104 10452 6132 10492
rect 6641 10489 6653 10492
rect 6687 10489 6699 10523
rect 6641 10483 6699 10489
rect 7098 10480 7104 10532
rect 7156 10520 7162 10532
rect 11256 10520 11284 10560
rect 12066 10548 12072 10600
rect 12124 10588 12130 10600
rect 12802 10588 12808 10600
rect 12124 10560 12808 10588
rect 12124 10548 12130 10560
rect 12802 10548 12808 10560
rect 12860 10588 12866 10600
rect 13173 10591 13231 10597
rect 13173 10588 13185 10591
rect 12860 10560 13185 10588
rect 12860 10548 12866 10560
rect 13173 10557 13185 10560
rect 13219 10557 13231 10591
rect 13173 10551 13231 10557
rect 13538 10548 13544 10600
rect 13596 10548 13602 10600
rect 13924 10588 13952 10619
rect 13998 10616 14004 10668
rect 14056 10616 14062 10668
rect 14093 10659 14151 10665
rect 14093 10625 14105 10659
rect 14139 10656 14151 10659
rect 14182 10656 14188 10668
rect 14139 10628 14188 10656
rect 14139 10625 14151 10628
rect 14093 10619 14151 10625
rect 14182 10616 14188 10628
rect 14240 10616 14246 10668
rect 14292 10665 14320 10696
rect 14277 10659 14335 10665
rect 14277 10625 14289 10659
rect 14323 10625 14335 10659
rect 14384 10656 14412 10764
rect 15102 10752 15108 10804
rect 15160 10792 15166 10804
rect 15289 10795 15347 10801
rect 15289 10792 15301 10795
rect 15160 10764 15301 10792
rect 15160 10752 15166 10764
rect 15289 10761 15301 10764
rect 15335 10761 15347 10795
rect 15289 10755 15347 10761
rect 15470 10752 15476 10804
rect 15528 10792 15534 10804
rect 15528 10764 15608 10792
rect 15528 10752 15534 10764
rect 14826 10684 14832 10736
rect 14884 10724 14890 10736
rect 15580 10724 15608 10764
rect 15654 10752 15660 10804
rect 15712 10792 15718 10804
rect 17655 10795 17713 10801
rect 17655 10792 17667 10795
rect 15712 10764 17667 10792
rect 15712 10752 15718 10764
rect 17655 10761 17667 10764
rect 17701 10761 17713 10795
rect 17655 10755 17713 10761
rect 17770 10752 17776 10804
rect 17828 10792 17834 10804
rect 18414 10792 18420 10804
rect 17828 10764 18420 10792
rect 17828 10752 17834 10764
rect 18414 10752 18420 10764
rect 18472 10752 18478 10804
rect 16942 10724 16948 10736
rect 14884 10696 15424 10724
rect 15580 10696 16436 10724
rect 14884 10684 14890 10696
rect 15013 10659 15071 10665
rect 15013 10656 15025 10659
rect 14384 10628 15025 10656
rect 14277 10619 14335 10625
rect 15013 10625 15025 10628
rect 15059 10625 15071 10659
rect 15013 10619 15071 10625
rect 15102 10616 15108 10668
rect 15160 10616 15166 10668
rect 15396 10665 15424 10696
rect 15387 10659 15445 10665
rect 15387 10625 15399 10659
rect 15433 10625 15445 10659
rect 15387 10619 15445 10625
rect 15562 10616 15568 10668
rect 15620 10656 15626 10668
rect 16117 10659 16175 10665
rect 16117 10656 16129 10659
rect 15620 10628 16129 10656
rect 15620 10616 15626 10628
rect 16117 10625 16129 10628
rect 16163 10625 16175 10659
rect 16117 10619 16175 10625
rect 16206 10616 16212 10668
rect 16264 10656 16270 10668
rect 16408 10665 16436 10696
rect 16776 10696 16948 10724
rect 16776 10665 16804 10696
rect 16942 10684 16948 10696
rect 17000 10684 17006 10736
rect 17865 10727 17923 10733
rect 17865 10693 17877 10727
rect 17911 10693 17923 10727
rect 17865 10687 17923 10693
rect 16301 10659 16359 10665
rect 16301 10656 16313 10659
rect 16264 10628 16313 10656
rect 16264 10616 16270 10628
rect 16301 10625 16313 10628
rect 16347 10625 16359 10659
rect 16301 10619 16359 10625
rect 16393 10659 16451 10665
rect 16393 10625 16405 10659
rect 16439 10625 16451 10659
rect 16393 10619 16451 10625
rect 16761 10659 16819 10665
rect 16761 10625 16773 10659
rect 16807 10625 16819 10659
rect 17494 10656 17500 10668
rect 16761 10619 16819 10625
rect 16868 10628 17500 10656
rect 14458 10588 14464 10600
rect 13924 10560 14464 10588
rect 14458 10548 14464 10560
rect 14516 10548 14522 10600
rect 14645 10591 14703 10597
rect 14645 10557 14657 10591
rect 14691 10588 14703 10591
rect 14826 10588 14832 10600
rect 14691 10560 14832 10588
rect 14691 10557 14703 10560
rect 14645 10551 14703 10557
rect 14826 10548 14832 10560
rect 14884 10548 14890 10600
rect 15473 10591 15531 10597
rect 15473 10588 15485 10591
rect 14936 10560 15485 10588
rect 7156 10492 11284 10520
rect 7156 10480 7162 10492
rect 11514 10480 11520 10532
rect 11572 10520 11578 10532
rect 11609 10523 11667 10529
rect 11609 10520 11621 10523
rect 11572 10492 11621 10520
rect 11572 10480 11578 10492
rect 11609 10489 11621 10492
rect 11655 10489 11667 10523
rect 11609 10483 11667 10489
rect 11790 10480 11796 10532
rect 11848 10520 11854 10532
rect 13998 10520 14004 10532
rect 11848 10492 14004 10520
rect 11848 10480 11854 10492
rect 13998 10480 14004 10492
rect 14056 10480 14062 10532
rect 14550 10480 14556 10532
rect 14608 10520 14614 10532
rect 14936 10520 14964 10560
rect 15473 10557 15485 10560
rect 15519 10557 15531 10591
rect 16408 10588 16436 10619
rect 16868 10588 16896 10628
rect 17494 10616 17500 10628
rect 17552 10616 17558 10668
rect 17880 10656 17908 10687
rect 17954 10684 17960 10736
rect 18012 10684 18018 10736
rect 18046 10656 18052 10668
rect 17880 10628 18052 10656
rect 18046 10616 18052 10628
rect 18104 10616 18110 10668
rect 18325 10659 18383 10665
rect 18325 10625 18337 10659
rect 18371 10656 18383 10659
rect 19150 10656 19156 10668
rect 18371 10628 19156 10656
rect 18371 10625 18383 10628
rect 18325 10619 18383 10625
rect 19150 10616 19156 10628
rect 19208 10616 19214 10668
rect 16408 10560 16896 10588
rect 15473 10551 15531 10557
rect 17034 10548 17040 10600
rect 17092 10588 17098 10600
rect 18141 10591 18199 10597
rect 18141 10588 18153 10591
rect 17092 10560 18153 10588
rect 17092 10548 17098 10560
rect 18141 10557 18153 10560
rect 18187 10557 18199 10591
rect 18141 10551 18199 10557
rect 15749 10523 15807 10529
rect 15749 10520 15761 10523
rect 14608 10492 14964 10520
rect 15166 10492 15761 10520
rect 14608 10480 14614 10492
rect 5776 10424 6132 10452
rect 5776 10412 5782 10424
rect 6454 10412 6460 10464
rect 6512 10412 6518 10464
rect 6546 10412 6552 10464
rect 6604 10452 6610 10464
rect 7650 10452 7656 10464
rect 6604 10424 7656 10452
rect 6604 10412 6610 10424
rect 7650 10412 7656 10424
rect 7708 10412 7714 10464
rect 8018 10412 8024 10464
rect 8076 10452 8082 10464
rect 8294 10452 8300 10464
rect 8076 10424 8300 10452
rect 8076 10412 8082 10424
rect 8294 10412 8300 10424
rect 8352 10452 8358 10464
rect 10778 10452 10784 10464
rect 8352 10424 10784 10452
rect 8352 10412 8358 10424
rect 10778 10412 10784 10424
rect 10836 10412 10842 10464
rect 10962 10412 10968 10464
rect 11020 10452 11026 10464
rect 13262 10452 13268 10464
rect 11020 10424 13268 10452
rect 11020 10412 11026 10424
rect 13262 10412 13268 10424
rect 13320 10412 13326 10464
rect 13906 10412 13912 10464
rect 13964 10452 13970 10464
rect 15166 10452 15194 10492
rect 15749 10489 15761 10492
rect 15795 10489 15807 10523
rect 15749 10483 15807 10489
rect 17494 10480 17500 10532
rect 17552 10480 17558 10532
rect 13964 10424 15194 10452
rect 13964 10412 13970 10424
rect 15378 10412 15384 10464
rect 15436 10412 15442 10464
rect 15838 10412 15844 10464
rect 15896 10452 15902 10464
rect 15933 10455 15991 10461
rect 15933 10452 15945 10455
rect 15896 10424 15945 10452
rect 15896 10412 15902 10424
rect 15933 10421 15945 10424
rect 15979 10421 15991 10455
rect 15933 10415 15991 10421
rect 16298 10412 16304 10464
rect 16356 10452 16362 10464
rect 16853 10455 16911 10461
rect 16853 10452 16865 10455
rect 16356 10424 16865 10452
rect 16356 10412 16362 10424
rect 16853 10421 16865 10424
rect 16899 10421 16911 10455
rect 16853 10415 16911 10421
rect 17034 10412 17040 10464
rect 17092 10452 17098 10464
rect 17221 10455 17279 10461
rect 17221 10452 17233 10455
rect 17092 10424 17233 10452
rect 17092 10412 17098 10424
rect 17221 10421 17233 10424
rect 17267 10421 17279 10455
rect 17221 10415 17279 10421
rect 17681 10455 17739 10461
rect 17681 10421 17693 10455
rect 17727 10452 17739 10455
rect 17862 10452 17868 10464
rect 17727 10424 17868 10452
rect 17727 10421 17739 10424
rect 17681 10415 17739 10421
rect 17862 10412 17868 10424
rect 17920 10412 17926 10464
rect 18049 10455 18107 10461
rect 18049 10421 18061 10455
rect 18095 10452 18107 10455
rect 18138 10452 18144 10464
rect 18095 10424 18144 10452
rect 18095 10421 18107 10424
rect 18049 10415 18107 10421
rect 18138 10412 18144 10424
rect 18196 10412 18202 10464
rect 1104 10362 18860 10384
rect 1104 10310 1950 10362
rect 2002 10310 2014 10362
rect 2066 10310 2078 10362
rect 2130 10310 2142 10362
rect 2194 10310 2206 10362
rect 2258 10310 6950 10362
rect 7002 10310 7014 10362
rect 7066 10310 7078 10362
rect 7130 10310 7142 10362
rect 7194 10310 7206 10362
rect 7258 10310 11950 10362
rect 12002 10310 12014 10362
rect 12066 10310 12078 10362
rect 12130 10310 12142 10362
rect 12194 10310 12206 10362
rect 12258 10310 16950 10362
rect 17002 10310 17014 10362
rect 17066 10310 17078 10362
rect 17130 10310 17142 10362
rect 17194 10310 17206 10362
rect 17258 10310 18860 10362
rect 1104 10288 18860 10310
rect 1394 10208 1400 10260
rect 1452 10248 1458 10260
rect 1946 10248 1952 10260
rect 1452 10220 1952 10248
rect 1452 10208 1458 10220
rect 1946 10208 1952 10220
rect 2004 10208 2010 10260
rect 3970 10208 3976 10260
rect 4028 10248 4034 10260
rect 4065 10251 4123 10257
rect 4065 10248 4077 10251
rect 4028 10220 4077 10248
rect 4028 10208 4034 10220
rect 4065 10217 4077 10220
rect 4111 10217 4123 10251
rect 4065 10211 4123 10217
rect 4338 10208 4344 10260
rect 4396 10248 4402 10260
rect 4982 10248 4988 10260
rect 4396 10220 4988 10248
rect 4396 10208 4402 10220
rect 4982 10208 4988 10220
rect 5040 10208 5046 10260
rect 5092 10220 8156 10248
rect 1854 10140 1860 10192
rect 1912 10180 1918 10192
rect 2130 10180 2136 10192
rect 1912 10152 2136 10180
rect 1912 10140 1918 10152
rect 2130 10140 2136 10152
rect 2188 10140 2194 10192
rect 2222 10140 2228 10192
rect 2280 10180 2286 10192
rect 2590 10180 2596 10192
rect 2280 10152 2596 10180
rect 2280 10140 2286 10152
rect 2590 10140 2596 10152
rect 2648 10140 2654 10192
rect 3344 10152 3832 10180
rect 1670 10072 1676 10124
rect 1728 10112 1734 10124
rect 1949 10115 2007 10121
rect 1949 10112 1961 10115
rect 1728 10084 1961 10112
rect 1728 10072 1734 10084
rect 1949 10081 1961 10084
rect 1995 10081 2007 10115
rect 2866 10112 2872 10124
rect 1949 10075 2007 10081
rect 2792 10084 2872 10112
rect 1210 10004 1216 10056
rect 1268 10044 1274 10056
rect 1394 10044 1400 10056
rect 1268 10016 1400 10044
rect 1268 10004 1274 10016
rect 1394 10004 1400 10016
rect 1452 10004 1458 10056
rect 2792 10053 2820 10084
rect 2866 10072 2872 10084
rect 2924 10072 2930 10124
rect 2777 10047 2835 10053
rect 2777 10013 2789 10047
rect 2823 10013 2835 10047
rect 2777 10007 2835 10013
rect 3050 10004 3056 10056
rect 3108 10004 3114 10056
rect 3344 10053 3372 10152
rect 3804 10112 3832 10152
rect 3878 10140 3884 10192
rect 3936 10180 3942 10192
rect 5092 10180 5120 10220
rect 3936 10152 5120 10180
rect 3936 10140 3942 10152
rect 5350 10140 5356 10192
rect 5408 10180 5414 10192
rect 7101 10183 7159 10189
rect 7101 10180 7113 10183
rect 5408 10152 7113 10180
rect 5408 10140 5414 10152
rect 7101 10149 7113 10152
rect 7147 10149 7159 10183
rect 7742 10180 7748 10192
rect 7101 10143 7159 10149
rect 7208 10152 7748 10180
rect 6362 10112 6368 10124
rect 3804 10084 6368 10112
rect 6362 10072 6368 10084
rect 6420 10072 6426 10124
rect 7006 10112 7012 10124
rect 6472 10084 7012 10112
rect 3329 10047 3387 10053
rect 3329 10013 3341 10047
rect 3375 10013 3387 10047
rect 3329 10007 3387 10013
rect 3513 10047 3571 10053
rect 3513 10013 3525 10047
rect 3559 10013 3571 10047
rect 3513 10007 3571 10013
rect 2682 9936 2688 9988
rect 2740 9976 2746 9988
rect 3421 9979 3479 9985
rect 3421 9976 3433 9979
rect 2740 9948 3433 9976
rect 2740 9936 2746 9948
rect 3421 9945 3433 9948
rect 3467 9945 3479 9979
rect 3528 9976 3556 10007
rect 3602 10004 3608 10056
rect 3660 10044 3666 10056
rect 3973 10047 4031 10053
rect 3973 10044 3985 10047
rect 3660 10016 3985 10044
rect 3660 10004 3666 10016
rect 3973 10013 3985 10016
rect 4019 10013 4031 10047
rect 3973 10007 4031 10013
rect 4246 10004 4252 10056
rect 4304 10004 4310 10056
rect 5166 10004 5172 10056
rect 5224 10044 5230 10056
rect 6472 10044 6500 10084
rect 7006 10072 7012 10084
rect 7064 10072 7070 10124
rect 7208 10112 7236 10152
rect 7742 10140 7748 10152
rect 7800 10140 7806 10192
rect 8128 10180 8156 10220
rect 8202 10208 8208 10260
rect 8260 10248 8266 10260
rect 11514 10248 11520 10260
rect 8260 10220 11520 10248
rect 8260 10208 8266 10220
rect 11514 10208 11520 10220
rect 11572 10208 11578 10260
rect 12526 10208 12532 10260
rect 12584 10248 12590 10260
rect 12986 10248 12992 10260
rect 12584 10220 12992 10248
rect 12584 10208 12590 10220
rect 12986 10208 12992 10220
rect 13044 10208 13050 10260
rect 13262 10208 13268 10260
rect 13320 10248 13326 10260
rect 14182 10248 14188 10260
rect 13320 10220 14188 10248
rect 13320 10208 13326 10220
rect 14182 10208 14188 10220
rect 14240 10248 14246 10260
rect 15378 10248 15384 10260
rect 14240 10220 15384 10248
rect 14240 10208 14246 10220
rect 15378 10208 15384 10220
rect 15436 10208 15442 10260
rect 16114 10248 16120 10260
rect 15856 10220 16120 10248
rect 15856 10192 15884 10220
rect 16114 10208 16120 10220
rect 16172 10208 16178 10260
rect 16482 10248 16488 10260
rect 16292 10220 16488 10248
rect 15102 10180 15108 10192
rect 8128 10152 15108 10180
rect 15102 10140 15108 10152
rect 15160 10140 15166 10192
rect 15838 10140 15844 10192
rect 15896 10140 15902 10192
rect 16025 10183 16083 10189
rect 16025 10149 16037 10183
rect 16071 10180 16083 10183
rect 16292 10180 16320 10220
rect 16482 10208 16488 10220
rect 16540 10208 16546 10260
rect 16758 10208 16764 10260
rect 16816 10248 16822 10260
rect 16942 10248 16948 10260
rect 16816 10220 16948 10248
rect 16816 10208 16822 10220
rect 16942 10208 16948 10220
rect 17000 10208 17006 10260
rect 18141 10251 18199 10257
rect 18141 10217 18153 10251
rect 18187 10248 18199 10251
rect 18414 10248 18420 10260
rect 18187 10220 18420 10248
rect 18187 10217 18199 10220
rect 18141 10211 18199 10217
rect 18414 10208 18420 10220
rect 18472 10208 18478 10260
rect 19058 10180 19064 10192
rect 16071 10152 16320 10180
rect 16963 10152 17816 10180
rect 16071 10149 16083 10152
rect 16025 10143 16083 10149
rect 7116 10084 7236 10112
rect 7469 10115 7527 10121
rect 5224 10016 6500 10044
rect 5224 10004 5230 10016
rect 7116 9988 7144 10084
rect 7469 10081 7481 10115
rect 7515 10112 7527 10115
rect 7515 10084 9444 10112
rect 7515 10081 7527 10084
rect 7469 10075 7527 10081
rect 7668 10053 7788 10054
rect 7285 10047 7343 10053
rect 7285 10013 7297 10047
rect 7331 10013 7343 10047
rect 7285 10007 7343 10013
rect 7561 10047 7619 10053
rect 7561 10013 7573 10047
rect 7607 10013 7619 10047
rect 7561 10007 7619 10013
rect 7653 10047 7788 10053
rect 7653 10013 7665 10047
rect 7699 10026 7788 10047
rect 7699 10013 7711 10026
rect 7653 10007 7711 10013
rect 4982 9976 4988 9988
rect 3528 9948 3832 9976
rect 3421 9939 3479 9945
rect 1210 9868 1216 9920
rect 1268 9908 1274 9920
rect 3510 9908 3516 9920
rect 1268 9880 3516 9908
rect 1268 9868 1274 9880
rect 3510 9868 3516 9880
rect 3568 9868 3574 9920
rect 3804 9908 3832 9948
rect 4632 9948 4988 9976
rect 4632 9908 4660 9948
rect 4982 9936 4988 9948
rect 5040 9936 5046 9988
rect 5350 9936 5356 9988
rect 5408 9976 5414 9988
rect 5626 9976 5632 9988
rect 5408 9948 5632 9976
rect 5408 9936 5414 9948
rect 5626 9936 5632 9948
rect 5684 9936 5690 9988
rect 7098 9936 7104 9988
rect 7156 9936 7162 9988
rect 7300 9976 7328 10007
rect 7374 9976 7380 9988
rect 7300 9948 7380 9976
rect 7374 9936 7380 9948
rect 7432 9936 7438 9988
rect 3804 9880 4660 9908
rect 4706 9868 4712 9920
rect 4764 9908 4770 9920
rect 4890 9908 4896 9920
rect 4764 9880 4896 9908
rect 4764 9868 4770 9880
rect 4890 9868 4896 9880
rect 4948 9868 4954 9920
rect 5718 9868 5724 9920
rect 5776 9908 5782 9920
rect 6822 9908 6828 9920
rect 5776 9880 6828 9908
rect 5776 9868 5782 9880
rect 6822 9868 6828 9880
rect 6880 9868 6886 9920
rect 7576 9908 7604 10007
rect 7760 9976 7788 10026
rect 7849 10047 7907 10053
rect 7849 10013 7861 10047
rect 7895 10044 7907 10047
rect 8938 10044 8944 10056
rect 7895 10016 8944 10044
rect 7895 10013 7907 10016
rect 7849 10007 7907 10013
rect 8938 10004 8944 10016
rect 8996 10004 9002 10056
rect 9416 10044 9444 10084
rect 9490 10072 9496 10124
rect 9548 10112 9554 10124
rect 9548 10084 16146 10112
rect 9548 10072 9554 10084
rect 10042 10044 10048 10056
rect 9416 10016 10048 10044
rect 10042 10004 10048 10016
rect 10100 10004 10106 10056
rect 15102 10004 15108 10056
rect 15160 10044 15166 10056
rect 15286 10044 15292 10056
rect 15160 10016 15292 10044
rect 15160 10004 15166 10016
rect 15286 10004 15292 10016
rect 15344 10004 15350 10056
rect 16393 10047 16451 10053
rect 16393 10013 16405 10047
rect 16439 10044 16451 10047
rect 16482 10044 16488 10056
rect 16439 10016 16488 10044
rect 16439 10013 16451 10016
rect 16393 10007 16451 10013
rect 16482 10004 16488 10016
rect 16540 10004 16546 10056
rect 16963 10044 16991 10152
rect 17405 10115 17463 10121
rect 17405 10081 17417 10115
rect 17451 10112 17463 10115
rect 17678 10112 17684 10124
rect 17451 10084 17684 10112
rect 17451 10081 17463 10084
rect 17405 10075 17463 10081
rect 17678 10072 17684 10084
rect 17736 10072 17742 10124
rect 16592 10016 16991 10044
rect 7760 9948 7880 9976
rect 7638 9908 7644 9920
rect 7576 9880 7644 9908
rect 7638 9868 7644 9880
rect 7696 9868 7702 9920
rect 7852 9908 7880 9948
rect 9490 9936 9496 9988
rect 9548 9976 9554 9988
rect 13262 9976 13268 9988
rect 9548 9948 13268 9976
rect 9548 9936 9554 9948
rect 13262 9936 13268 9948
rect 13320 9936 13326 9988
rect 15378 9936 15384 9988
rect 15436 9976 15442 9988
rect 16592 9976 16620 10016
rect 17034 10004 17040 10056
rect 17092 10004 17098 10056
rect 17494 10004 17500 10056
rect 17552 10004 17558 10056
rect 17589 10047 17647 10053
rect 17589 10013 17601 10047
rect 17635 10013 17647 10047
rect 17589 10007 17647 10013
rect 15436 9948 16620 9976
rect 15436 9936 15442 9948
rect 16666 9936 16672 9988
rect 16724 9976 16730 9988
rect 17604 9976 17632 10007
rect 16724 9948 17632 9976
rect 16724 9936 16730 9948
rect 8938 9908 8944 9920
rect 7852 9880 8944 9908
rect 8938 9868 8944 9880
rect 8996 9868 9002 9920
rect 12342 9868 12348 9920
rect 12400 9908 12406 9920
rect 12618 9908 12624 9920
rect 12400 9880 12624 9908
rect 12400 9868 12406 9880
rect 12618 9868 12624 9880
rect 12676 9868 12682 9920
rect 12802 9868 12808 9920
rect 12860 9908 12866 9920
rect 14826 9908 14832 9920
rect 12860 9880 14832 9908
rect 12860 9868 12866 9880
rect 14826 9868 14832 9880
rect 14884 9868 14890 9920
rect 17494 9868 17500 9920
rect 17552 9908 17558 9920
rect 17696 9908 17724 10072
rect 17788 10044 17816 10152
rect 17972 10152 19064 10180
rect 17972 10053 18000 10152
rect 19058 10140 19064 10152
rect 19116 10140 19122 10192
rect 18138 10072 18144 10124
rect 18196 10112 18202 10124
rect 18305 10115 18363 10121
rect 18305 10112 18317 10115
rect 18196 10084 18317 10112
rect 18196 10072 18202 10084
rect 18305 10081 18317 10084
rect 18351 10081 18363 10115
rect 18305 10075 18363 10081
rect 17865 10047 17923 10053
rect 17865 10044 17877 10047
rect 17788 10016 17877 10044
rect 17865 10013 17877 10016
rect 17911 10013 17923 10047
rect 17865 10007 17923 10013
rect 17957 10047 18015 10053
rect 17957 10013 17969 10047
rect 18003 10013 18015 10047
rect 18509 10047 18567 10053
rect 18509 10044 18521 10047
rect 17957 10007 18015 10013
rect 18064 10016 18521 10044
rect 17770 9936 17776 9988
rect 17828 9936 17834 9988
rect 17880 9976 17908 10007
rect 18064 9976 18092 10016
rect 18509 10013 18521 10016
rect 18555 10013 18567 10047
rect 18509 10007 18567 10013
rect 17880 9948 18092 9976
rect 18233 9979 18291 9985
rect 18233 9945 18245 9979
rect 18279 9976 18291 9979
rect 18874 9976 18880 9988
rect 18279 9948 18880 9976
rect 18279 9945 18291 9948
rect 18233 9939 18291 9945
rect 18874 9936 18880 9948
rect 18932 9936 18938 9988
rect 17552 9880 17724 9908
rect 17788 9908 17816 9936
rect 18417 9911 18475 9917
rect 18417 9908 18429 9911
rect 17788 9880 18429 9908
rect 17552 9868 17558 9880
rect 18417 9877 18429 9880
rect 18463 9877 18475 9911
rect 18417 9871 18475 9877
rect 1104 9818 18860 9840
rect 1104 9766 2610 9818
rect 2662 9766 2674 9818
rect 2726 9766 2738 9818
rect 2790 9766 2802 9818
rect 2854 9766 2866 9818
rect 2918 9766 7610 9818
rect 7662 9766 7674 9818
rect 7726 9766 7738 9818
rect 7790 9766 7802 9818
rect 7854 9766 7866 9818
rect 7918 9766 12610 9818
rect 12662 9766 12674 9818
rect 12726 9766 12738 9818
rect 12790 9766 12802 9818
rect 12854 9766 12866 9818
rect 12918 9766 17610 9818
rect 17662 9766 17674 9818
rect 17726 9766 17738 9818
rect 17790 9766 17802 9818
rect 17854 9766 17866 9818
rect 17918 9766 18860 9818
rect 1104 9744 18860 9766
rect 106 9664 112 9716
rect 164 9704 170 9716
rect 164 9676 2360 9704
rect 164 9664 170 9676
rect 1026 9596 1032 9648
rect 1084 9636 1090 9648
rect 1578 9636 1584 9648
rect 1084 9608 1584 9636
rect 1084 9596 1090 9608
rect 1578 9596 1584 9608
rect 1636 9596 1642 9648
rect 2332 9636 2360 9676
rect 2406 9664 2412 9716
rect 2464 9704 2470 9716
rect 2590 9704 2596 9716
rect 2464 9676 2596 9704
rect 2464 9664 2470 9676
rect 2590 9664 2596 9676
rect 2648 9664 2654 9716
rect 2700 9676 4200 9704
rect 2700 9636 2728 9676
rect 1688 9608 1900 9636
rect 2332 9608 2728 9636
rect 382 9528 388 9580
rect 440 9568 446 9580
rect 1688 9568 1716 9608
rect 1872 9577 1900 9608
rect 2866 9596 2872 9648
rect 2924 9596 2930 9648
rect 3786 9636 3792 9648
rect 2976 9608 3792 9636
rect 440 9540 1716 9568
rect 1765 9571 1823 9577
rect 440 9528 446 9540
rect 1765 9537 1777 9571
rect 1811 9537 1823 9571
rect 1765 9531 1823 9537
rect 1857 9571 1915 9577
rect 1857 9537 1869 9571
rect 1903 9537 1915 9571
rect 1857 9531 1915 9537
rect 1780 9500 1808 9531
rect 2038 9528 2044 9580
rect 2096 9528 2102 9580
rect 2406 9528 2412 9580
rect 2464 9568 2470 9580
rect 2501 9571 2559 9577
rect 2501 9568 2513 9571
rect 2464 9540 2513 9568
rect 2464 9528 2470 9540
rect 2501 9537 2513 9540
rect 2547 9537 2559 9571
rect 2774 9568 2780 9580
rect 2501 9531 2559 9537
rect 2608 9540 2780 9568
rect 2608 9500 2636 9540
rect 2774 9528 2780 9540
rect 2832 9568 2838 9580
rect 2976 9568 3004 9608
rect 3786 9596 3792 9608
rect 3844 9596 3850 9648
rect 4172 9636 4200 9676
rect 4246 9664 4252 9716
rect 4304 9704 4310 9716
rect 4304 9676 5764 9704
rect 4304 9664 4310 9676
rect 4801 9639 4859 9645
rect 4801 9636 4813 9639
rect 4172 9608 4813 9636
rect 4801 9605 4813 9608
rect 4847 9605 4859 9639
rect 4801 9599 4859 9605
rect 2832 9540 3004 9568
rect 2832 9528 2838 9540
rect 3050 9528 3056 9580
rect 3108 9528 3114 9580
rect 3878 9568 3884 9580
rect 3160 9540 3884 9568
rect 1780 9472 2636 9500
rect 2866 9460 2872 9512
rect 2924 9500 2930 9512
rect 3160 9500 3188 9540
rect 3878 9528 3884 9540
rect 3936 9528 3942 9580
rect 4617 9571 4675 9577
rect 4617 9537 4629 9571
rect 4663 9537 4675 9571
rect 4617 9531 4675 9537
rect 4893 9571 4951 9577
rect 4893 9537 4905 9571
rect 4939 9568 4951 9571
rect 5626 9568 5632 9580
rect 4939 9540 5632 9568
rect 4939 9537 4951 9540
rect 4893 9531 4951 9537
rect 2924 9472 3188 9500
rect 2924 9460 2930 9472
rect 3326 9460 3332 9512
rect 3384 9460 3390 9512
rect 3510 9460 3516 9512
rect 3568 9500 3574 9512
rect 3789 9503 3847 9509
rect 3789 9500 3801 9503
rect 3568 9472 3801 9500
rect 3568 9460 3574 9472
rect 3789 9469 3801 9472
rect 3835 9500 3847 9503
rect 4246 9500 4252 9512
rect 3835 9472 4252 9500
rect 3835 9469 3847 9472
rect 3789 9463 3847 9469
rect 4246 9460 4252 9472
rect 4304 9500 4310 9512
rect 4433 9503 4491 9509
rect 4433 9500 4445 9503
rect 4304 9472 4445 9500
rect 4304 9460 4310 9472
rect 4433 9469 4445 9472
rect 4479 9469 4491 9503
rect 4632 9500 4660 9531
rect 5626 9528 5632 9540
rect 5684 9528 5690 9580
rect 5736 9568 5764 9676
rect 5902 9664 5908 9716
rect 5960 9704 5966 9716
rect 6178 9704 6184 9716
rect 5960 9676 6184 9704
rect 5960 9664 5966 9676
rect 6178 9664 6184 9676
rect 6236 9664 6242 9716
rect 6362 9664 6368 9716
rect 6420 9704 6426 9716
rect 9030 9704 9036 9716
rect 6420 9676 9036 9704
rect 6420 9664 6426 9676
rect 9030 9664 9036 9676
rect 9088 9704 9094 9716
rect 10962 9704 10968 9716
rect 9088 9676 10968 9704
rect 9088 9664 9094 9676
rect 10962 9664 10968 9676
rect 11020 9664 11026 9716
rect 11054 9664 11060 9716
rect 11112 9704 11118 9716
rect 12158 9704 12164 9716
rect 11112 9676 12164 9704
rect 11112 9664 11118 9676
rect 12158 9664 12164 9676
rect 12216 9664 12222 9716
rect 12250 9664 12256 9716
rect 12308 9664 12314 9716
rect 13262 9664 13268 9716
rect 13320 9704 13326 9716
rect 15102 9704 15108 9716
rect 13320 9676 15108 9704
rect 13320 9664 13326 9676
rect 15102 9664 15108 9676
rect 15160 9704 15166 9716
rect 17218 9704 17224 9716
rect 15160 9676 17224 9704
rect 15160 9664 15166 9676
rect 17218 9664 17224 9676
rect 17276 9664 17282 9716
rect 6822 9636 6828 9648
rect 5920 9608 6828 9636
rect 5920 9568 5948 9608
rect 6822 9596 6828 9608
rect 6880 9596 6886 9648
rect 12342 9636 12348 9648
rect 7392 9608 9076 9636
rect 7392 9602 7420 9608
rect 5736 9540 5948 9568
rect 6178 9528 6184 9580
rect 6236 9568 6242 9580
rect 7098 9568 7104 9580
rect 6236 9540 7104 9568
rect 6236 9528 6242 9540
rect 7098 9528 7104 9540
rect 7156 9528 7162 9580
rect 7208 9577 7420 9602
rect 9048 9580 9076 9608
rect 10520 9608 12348 9636
rect 7193 9574 7420 9577
rect 7193 9571 7251 9574
rect 7193 9537 7205 9571
rect 7239 9537 7251 9571
rect 7193 9531 7251 9537
rect 5166 9500 5172 9512
rect 4632 9472 5172 9500
rect 4433 9463 4491 9469
rect 5166 9460 5172 9472
rect 5224 9460 5230 9512
rect 6362 9460 6368 9512
rect 6420 9500 6426 9512
rect 7208 9500 7236 9531
rect 7742 9528 7748 9580
rect 7800 9528 7806 9580
rect 9030 9528 9036 9580
rect 9088 9528 9094 9580
rect 9490 9528 9496 9580
rect 9548 9568 9554 9580
rect 9585 9571 9643 9577
rect 9585 9568 9597 9571
rect 9548 9540 9597 9568
rect 9548 9528 9554 9540
rect 9585 9537 9597 9540
rect 9631 9537 9643 9571
rect 9585 9531 9643 9537
rect 9953 9571 10011 9577
rect 9953 9537 9965 9571
rect 9999 9537 10011 9571
rect 9953 9531 10011 9537
rect 6420 9472 7236 9500
rect 7561 9503 7619 9509
rect 6420 9460 6426 9472
rect 7561 9469 7573 9503
rect 7607 9500 7619 9503
rect 7650 9500 7656 9512
rect 7607 9472 7656 9500
rect 7607 9469 7619 9472
rect 7561 9463 7619 9469
rect 7650 9460 7656 9472
rect 7708 9460 7714 9512
rect 7926 9460 7932 9512
rect 7984 9500 7990 9512
rect 8941 9503 8999 9509
rect 8941 9500 8953 9503
rect 7984 9472 8953 9500
rect 7984 9460 7990 9472
rect 8941 9469 8953 9472
rect 8987 9469 8999 9503
rect 8941 9463 8999 9469
rect 9677 9503 9735 9509
rect 9677 9469 9689 9503
rect 9723 9500 9735 9503
rect 9766 9500 9772 9512
rect 9723 9472 9772 9500
rect 9723 9469 9735 9472
rect 9677 9463 9735 9469
rect 9766 9460 9772 9472
rect 9824 9460 9830 9512
rect 9861 9503 9919 9509
rect 9861 9469 9873 9503
rect 9907 9469 9919 9503
rect 9968 9500 9996 9531
rect 10318 9528 10324 9580
rect 10376 9528 10382 9580
rect 10520 9500 10548 9608
rect 12342 9596 12348 9608
rect 12400 9636 12406 9648
rect 12802 9636 12808 9648
rect 12400 9608 12808 9636
rect 12400 9596 12406 9608
rect 12802 9596 12808 9608
rect 12860 9596 12866 9648
rect 14829 9639 14887 9645
rect 14829 9605 14841 9639
rect 14875 9636 14887 9639
rect 14875 9608 15148 9636
rect 14875 9605 14887 9608
rect 14829 9599 14887 9605
rect 10594 9528 10600 9580
rect 10652 9568 10658 9580
rect 10778 9568 10784 9580
rect 10652 9540 10784 9568
rect 10652 9528 10658 9540
rect 10778 9528 10784 9540
rect 10836 9568 10842 9580
rect 12161 9571 12219 9577
rect 12161 9568 12173 9571
rect 10836 9540 12173 9568
rect 10836 9528 10842 9540
rect 12161 9537 12173 9540
rect 12207 9537 12219 9571
rect 12161 9531 12219 9537
rect 12526 9528 12532 9580
rect 12584 9568 12590 9580
rect 13909 9571 13967 9577
rect 13909 9568 13921 9571
rect 12584 9540 13921 9568
rect 12584 9528 12590 9540
rect 13909 9537 13921 9540
rect 13955 9537 13967 9571
rect 13909 9531 13967 9537
rect 14001 9571 14059 9577
rect 14001 9537 14013 9571
rect 14047 9537 14059 9571
rect 14001 9531 14059 9537
rect 14182 9534 14188 9586
rect 14240 9534 14246 9586
rect 15120 9580 15148 9608
rect 16942 9596 16948 9648
rect 17000 9596 17006 9648
rect 17402 9636 17408 9648
rect 17144 9608 17408 9636
rect 14458 9568 14464 9580
rect 14292 9540 14464 9568
rect 14185 9531 14243 9534
rect 9968 9472 10548 9500
rect 9861 9463 9919 9469
rect 2130 9392 2136 9444
rect 2188 9432 2194 9444
rect 3237 9435 3295 9441
rect 2188 9404 3188 9432
rect 2188 9392 2194 9404
rect 1670 9324 1676 9376
rect 1728 9364 1734 9376
rect 2041 9367 2099 9373
rect 2041 9364 2053 9367
rect 1728 9336 2053 9364
rect 1728 9324 1734 9336
rect 2041 9333 2053 9336
rect 2087 9364 2099 9367
rect 2222 9364 2228 9376
rect 2087 9336 2228 9364
rect 2087 9333 2099 9336
rect 2041 9327 2099 9333
rect 2222 9324 2228 9336
rect 2280 9324 2286 9376
rect 2682 9324 2688 9376
rect 2740 9324 2746 9376
rect 3160 9364 3188 9404
rect 3237 9401 3249 9435
rect 3283 9432 3295 9435
rect 3283 9404 6040 9432
rect 3283 9401 3295 9404
rect 3237 9395 3295 9401
rect 3602 9364 3608 9376
rect 3160 9336 3608 9364
rect 3602 9324 3608 9336
rect 3660 9324 3666 9376
rect 4249 9367 4307 9373
rect 4249 9333 4261 9367
rect 4295 9364 4307 9367
rect 5166 9364 5172 9376
rect 4295 9336 5172 9364
rect 4295 9333 4307 9336
rect 4249 9327 4307 9333
rect 5166 9324 5172 9336
rect 5224 9324 5230 9376
rect 6012 9364 6040 9404
rect 6748 9404 9536 9432
rect 6748 9364 6776 9404
rect 6012 9336 6776 9364
rect 6822 9324 6828 9376
rect 6880 9364 6886 9376
rect 8202 9364 8208 9376
rect 6880 9336 8208 9364
rect 6880 9324 6886 9336
rect 8202 9324 8208 9336
rect 8260 9324 8266 9376
rect 9508 9364 9536 9404
rect 9582 9392 9588 9444
rect 9640 9432 9646 9444
rect 9876 9432 9904 9463
rect 10870 9460 10876 9512
rect 10928 9460 10934 9512
rect 11238 9460 11244 9512
rect 11296 9500 11302 9512
rect 14016 9500 14044 9531
rect 14292 9500 14320 9540
rect 14458 9528 14464 9540
rect 14516 9528 14522 9580
rect 14645 9571 14703 9577
rect 14645 9537 14657 9571
rect 14691 9537 14703 9571
rect 14645 9531 14703 9537
rect 11296 9472 14044 9500
rect 14117 9472 14320 9500
rect 14660 9500 14688 9531
rect 14734 9528 14740 9580
rect 14792 9568 14798 9580
rect 14921 9571 14979 9577
rect 14921 9568 14933 9571
rect 14792 9540 14933 9568
rect 14792 9528 14798 9540
rect 14921 9537 14933 9540
rect 14967 9537 14979 9571
rect 14921 9531 14979 9537
rect 15102 9528 15108 9580
rect 15160 9528 15166 9580
rect 15930 9528 15936 9580
rect 15988 9568 15994 9580
rect 15988 9540 16344 9568
rect 15988 9528 15994 9540
rect 15470 9500 15476 9512
rect 14660 9472 15476 9500
rect 11296 9460 11302 9472
rect 10888 9432 10916 9460
rect 9640 9404 10916 9432
rect 9640 9392 9646 9404
rect 10962 9392 10968 9444
rect 11020 9432 11026 9444
rect 12526 9432 12532 9444
rect 11020 9404 12532 9432
rect 11020 9392 11026 9404
rect 12526 9392 12532 9404
rect 12584 9392 12590 9444
rect 12986 9392 12992 9444
rect 13044 9432 13050 9444
rect 14117 9432 14145 9472
rect 15470 9460 15476 9472
rect 15528 9500 15534 9512
rect 16206 9500 16212 9512
rect 15528 9472 16212 9500
rect 15528 9460 15534 9472
rect 16206 9460 16212 9472
rect 16264 9460 16270 9512
rect 16316 9500 16344 9540
rect 16482 9528 16488 9580
rect 16540 9568 16546 9580
rect 16669 9571 16727 9577
rect 16669 9568 16681 9571
rect 16540 9540 16681 9568
rect 16540 9528 16546 9540
rect 16669 9537 16681 9540
rect 16715 9537 16727 9571
rect 16669 9531 16727 9537
rect 16780 9571 16838 9577
rect 16780 9537 16792 9571
rect 16826 9568 16838 9571
rect 17144 9568 17172 9608
rect 17402 9596 17408 9608
rect 17460 9596 17466 9648
rect 16826 9540 17172 9568
rect 16826 9537 16838 9540
rect 16780 9531 16838 9537
rect 17218 9528 17224 9580
rect 17276 9528 17282 9580
rect 17770 9528 17776 9580
rect 17828 9528 17834 9580
rect 18138 9528 18144 9580
rect 18196 9568 18202 9580
rect 19334 9568 19340 9580
rect 18196 9540 19340 9568
rect 18196 9528 18202 9540
rect 19334 9528 19340 9540
rect 19392 9528 19398 9580
rect 17405 9503 17463 9509
rect 17405 9500 17417 9503
rect 16316 9472 17417 9500
rect 13044 9404 14145 9432
rect 13044 9392 13050 9404
rect 14458 9392 14464 9444
rect 14516 9392 14522 9444
rect 15930 9432 15936 9444
rect 14660 9404 15936 9432
rect 10594 9364 10600 9376
rect 9508 9336 10600 9364
rect 10594 9324 10600 9336
rect 10652 9324 10658 9376
rect 10686 9324 10692 9376
rect 10744 9364 10750 9376
rect 11698 9364 11704 9376
rect 10744 9336 11704 9364
rect 10744 9324 10750 9336
rect 11698 9324 11704 9336
rect 11756 9324 11762 9376
rect 11882 9324 11888 9376
rect 11940 9364 11946 9376
rect 12342 9364 12348 9376
rect 11940 9336 12348 9364
rect 11940 9324 11946 9336
rect 12342 9324 12348 9336
rect 12400 9324 12406 9376
rect 14274 9324 14280 9376
rect 14332 9364 14338 9376
rect 14369 9367 14427 9373
rect 14369 9364 14381 9367
rect 14332 9336 14381 9364
rect 14332 9324 14338 9336
rect 14369 9333 14381 9336
rect 14415 9364 14427 9367
rect 14660 9364 14688 9404
rect 15930 9392 15936 9404
rect 15988 9392 15994 9444
rect 16316 9432 16344 9472
rect 17405 9469 17417 9472
rect 17451 9469 17463 9503
rect 17405 9463 17463 9469
rect 16040 9404 16344 9432
rect 14415 9336 14688 9364
rect 14415 9333 14427 9336
rect 14369 9327 14427 9333
rect 14734 9324 14740 9376
rect 14792 9364 14798 9376
rect 16040 9364 16068 9404
rect 16482 9392 16488 9444
rect 16540 9432 16546 9444
rect 16540 9404 16804 9432
rect 16540 9392 16546 9404
rect 14792 9336 16068 9364
rect 14792 9324 14798 9336
rect 16298 9324 16304 9376
rect 16356 9364 16362 9376
rect 16669 9367 16727 9373
rect 16669 9364 16681 9367
rect 16356 9336 16681 9364
rect 16356 9324 16362 9336
rect 16669 9333 16681 9336
rect 16715 9333 16727 9367
rect 16776 9364 16804 9404
rect 17770 9364 17776 9376
rect 16776 9336 17776 9364
rect 16669 9327 16727 9333
rect 17770 9324 17776 9336
rect 17828 9324 17834 9376
rect 1104 9274 18860 9296
rect 1104 9222 1950 9274
rect 2002 9222 2014 9274
rect 2066 9222 2078 9274
rect 2130 9222 2142 9274
rect 2194 9222 2206 9274
rect 2258 9222 6950 9274
rect 7002 9222 7014 9274
rect 7066 9222 7078 9274
rect 7130 9222 7142 9274
rect 7194 9222 7206 9274
rect 7258 9222 11950 9274
rect 12002 9222 12014 9274
rect 12066 9222 12078 9274
rect 12130 9222 12142 9274
rect 12194 9222 12206 9274
rect 12258 9222 16950 9274
rect 17002 9222 17014 9274
rect 17066 9222 17078 9274
rect 17130 9222 17142 9274
rect 17194 9222 17206 9274
rect 17258 9222 18860 9274
rect 1104 9200 18860 9222
rect 1397 9163 1455 9169
rect 1397 9129 1409 9163
rect 1443 9160 1455 9163
rect 2406 9160 2412 9172
rect 1443 9132 2412 9160
rect 1443 9129 1455 9132
rect 1397 9123 1455 9129
rect 2406 9120 2412 9132
rect 2464 9120 2470 9172
rect 2498 9120 2504 9172
rect 2556 9160 2562 9172
rect 2685 9163 2743 9169
rect 2685 9160 2697 9163
rect 2556 9132 2697 9160
rect 2556 9120 2562 9132
rect 2685 9129 2697 9132
rect 2731 9129 2743 9163
rect 3418 9160 3424 9172
rect 2685 9123 2743 9129
rect 2976 9132 3424 9160
rect 2976 9024 3004 9132
rect 3418 9120 3424 9132
rect 3476 9120 3482 9172
rect 3786 9120 3792 9172
rect 3844 9160 3850 9172
rect 4154 9160 4160 9172
rect 3844 9132 4160 9160
rect 3844 9120 3850 9132
rect 4154 9120 4160 9132
rect 4212 9120 4218 9172
rect 4816 9132 5028 9160
rect 3145 9095 3203 9101
rect 3145 9061 3157 9095
rect 3191 9092 3203 9095
rect 3191 9064 3832 9092
rect 3191 9061 3203 9064
rect 3145 9055 3203 9061
rect 3804 9024 3832 9064
rect 3878 9052 3884 9104
rect 3936 9092 3942 9104
rect 4816 9092 4844 9132
rect 3936 9064 4844 9092
rect 5000 9092 5028 9132
rect 5074 9120 5080 9172
rect 5132 9160 5138 9172
rect 6822 9160 6828 9172
rect 5132 9132 6828 9160
rect 5132 9120 5138 9132
rect 6822 9120 6828 9132
rect 6880 9120 6886 9172
rect 7742 9120 7748 9172
rect 7800 9160 7806 9172
rect 8386 9160 8392 9172
rect 7800 9132 8392 9160
rect 7800 9120 7806 9132
rect 8386 9120 8392 9132
rect 8444 9120 8450 9172
rect 9766 9120 9772 9172
rect 9824 9160 9830 9172
rect 10686 9160 10692 9172
rect 9824 9132 10692 9160
rect 9824 9120 9830 9132
rect 10686 9120 10692 9132
rect 10744 9120 10750 9172
rect 10965 9163 11023 9169
rect 10965 9129 10977 9163
rect 11011 9160 11023 9163
rect 11330 9160 11336 9172
rect 11011 9132 11336 9160
rect 11011 9129 11023 9132
rect 10965 9123 11023 9129
rect 11330 9120 11336 9132
rect 11388 9120 11394 9172
rect 11606 9120 11612 9172
rect 11664 9160 11670 9172
rect 12158 9160 12164 9172
rect 11664 9132 12164 9160
rect 11664 9120 11670 9132
rect 12158 9120 12164 9132
rect 12216 9120 12222 9172
rect 12434 9120 12440 9172
rect 12492 9160 12498 9172
rect 13630 9160 13636 9172
rect 12492 9132 13636 9160
rect 12492 9120 12498 9132
rect 13630 9120 13636 9132
rect 13688 9160 13694 9172
rect 14458 9160 14464 9172
rect 13688 9132 14464 9160
rect 13688 9120 13694 9132
rect 14458 9120 14464 9132
rect 14516 9120 14522 9172
rect 18230 9160 18236 9172
rect 14844 9132 18236 9160
rect 10781 9095 10839 9101
rect 10781 9092 10793 9095
rect 5000 9064 10793 9092
rect 3936 9052 3942 9064
rect 10781 9061 10793 9064
rect 10827 9061 10839 9095
rect 10781 9055 10839 9061
rect 10870 9052 10876 9104
rect 10928 9092 10934 9104
rect 13722 9092 13728 9104
rect 10928 9064 13728 9092
rect 10928 9052 10934 9064
rect 13722 9052 13728 9064
rect 13780 9052 13786 9104
rect 13906 9052 13912 9104
rect 13964 9092 13970 9104
rect 14844 9092 14872 9132
rect 18230 9120 18236 9132
rect 18288 9120 18294 9172
rect 13964 9064 14872 9092
rect 13964 9052 13970 9064
rect 14918 9052 14924 9104
rect 14976 9092 14982 9104
rect 15194 9092 15200 9104
rect 14976 9064 15200 9092
rect 14976 9052 14982 9064
rect 15194 9052 15200 9064
rect 15252 9052 15258 9104
rect 16758 9092 16764 9104
rect 16316 9064 16764 9092
rect 7098 9024 7104 9036
rect 2884 8996 3004 9024
rect 3344 8996 3648 9024
rect 3804 8996 7104 9024
rect 1578 8916 1584 8968
rect 1636 8916 1642 8968
rect 1857 8959 1915 8965
rect 1857 8925 1869 8959
rect 1903 8925 1915 8959
rect 1857 8919 1915 8925
rect 750 8848 756 8900
rect 808 8888 814 8900
rect 1872 8888 1900 8919
rect 1946 8916 1952 8968
rect 2004 8916 2010 8968
rect 2884 8965 2912 8996
rect 2869 8959 2927 8965
rect 2869 8925 2881 8959
rect 2915 8925 2927 8959
rect 2869 8919 2927 8925
rect 2958 8916 2964 8968
rect 3016 8916 3022 8968
rect 3344 8965 3372 8996
rect 3620 8966 3648 8996
rect 7098 8984 7104 8996
rect 7156 8984 7162 9036
rect 7374 8984 7380 9036
rect 7432 9024 7438 9036
rect 7432 8996 7696 9024
rect 7432 8984 7438 8996
rect 3237 8959 3295 8965
rect 3237 8925 3249 8959
rect 3283 8925 3295 8959
rect 3237 8919 3295 8925
rect 3329 8959 3387 8965
rect 3329 8925 3341 8959
rect 3375 8925 3387 8959
rect 3620 8956 3740 8966
rect 4062 8956 4068 8968
rect 3620 8938 4068 8956
rect 3712 8928 4068 8938
rect 3329 8919 3387 8925
rect 808 8860 1900 8888
rect 808 8848 814 8860
rect 2222 8848 2228 8900
rect 2280 8848 2286 8900
rect 2406 8848 2412 8900
rect 2464 8888 2470 8900
rect 3252 8888 3280 8919
rect 4062 8916 4068 8928
rect 4120 8916 4126 8968
rect 4154 8916 4160 8968
rect 4212 8916 4218 8968
rect 4246 8916 4252 8968
rect 4304 8956 4310 8968
rect 4433 8959 4491 8965
rect 4433 8956 4445 8959
rect 4304 8928 4445 8956
rect 4304 8916 4310 8928
rect 4433 8925 4445 8928
rect 4479 8925 4491 8959
rect 4433 8919 4491 8925
rect 4614 8916 4620 8968
rect 4672 8956 4678 8968
rect 4801 8959 4859 8965
rect 4801 8956 4813 8959
rect 4672 8928 4813 8956
rect 4672 8916 4678 8928
rect 4801 8925 4813 8928
rect 4847 8925 4859 8959
rect 4801 8919 4859 8925
rect 4893 8959 4951 8965
rect 4893 8925 4905 8959
rect 4939 8925 4951 8959
rect 4893 8919 4951 8925
rect 2464 8860 3280 8888
rect 3513 8891 3571 8897
rect 2464 8848 2470 8860
rect 3513 8857 3525 8891
rect 3559 8888 3571 8891
rect 3602 8888 3608 8900
rect 3559 8860 3608 8888
rect 3559 8857 3571 8860
rect 3513 8851 3571 8857
rect 3602 8848 3608 8860
rect 3660 8848 3666 8900
rect 3878 8848 3884 8900
rect 3936 8848 3942 8900
rect 4172 8888 4200 8916
rect 4172 8860 4292 8888
rect 4264 8832 4292 8860
rect 4908 8832 4936 8919
rect 5074 8916 5080 8968
rect 5132 8916 5138 8968
rect 5169 8959 5227 8965
rect 5169 8925 5181 8959
rect 5215 8950 5227 8959
rect 5258 8950 5264 8968
rect 5215 8925 5264 8950
rect 5169 8922 5264 8925
rect 5169 8919 5227 8922
rect 5258 8916 5264 8922
rect 5316 8916 5322 8968
rect 5350 8916 5356 8968
rect 5408 8916 5414 8968
rect 6362 8916 6368 8968
rect 6420 8956 6426 8968
rect 7561 8959 7619 8965
rect 7561 8956 7573 8959
rect 6420 8928 7573 8956
rect 6420 8916 6426 8928
rect 7561 8925 7573 8928
rect 7607 8925 7619 8959
rect 7668 8942 7696 8996
rect 8110 8984 8116 9036
rect 8168 9024 8174 9036
rect 8481 9027 8539 9033
rect 8481 9024 8493 9027
rect 8168 8996 8493 9024
rect 8168 8984 8174 8996
rect 8481 8993 8493 8996
rect 8527 9024 8539 9027
rect 8570 9024 8576 9036
rect 8527 8996 8576 9024
rect 8527 8993 8539 8996
rect 8481 8987 8539 8993
rect 8570 8984 8576 8996
rect 8628 8984 8634 9036
rect 9030 8984 9036 9036
rect 9088 9024 9094 9036
rect 9214 9024 9220 9036
rect 9088 8996 9220 9024
rect 9088 8984 9094 8996
rect 9214 8984 9220 8996
rect 9272 8984 9278 9036
rect 10318 9024 10324 9036
rect 10060 8996 10324 9024
rect 7561 8919 7619 8925
rect 5368 8888 5396 8916
rect 7926 8888 7932 8900
rect 5368 8860 7932 8888
rect 7926 8848 7932 8860
rect 7984 8848 7990 8900
rect 8110 8848 8116 8900
rect 8168 8888 8174 8900
rect 8941 8891 8999 8897
rect 8941 8888 8953 8891
rect 8168 8860 8953 8888
rect 8168 8848 8174 8860
rect 8941 8857 8953 8860
rect 8987 8888 8999 8891
rect 9950 8888 9956 8900
rect 8987 8860 9956 8888
rect 8987 8857 8999 8860
rect 8941 8851 8999 8857
rect 9950 8848 9956 8860
rect 10008 8848 10014 8900
rect 1118 8780 1124 8832
rect 1176 8820 1182 8832
rect 1578 8820 1584 8832
rect 1176 8792 1584 8820
rect 1176 8780 1182 8792
rect 1578 8780 1584 8792
rect 1636 8820 1642 8832
rect 1765 8823 1823 8829
rect 1765 8820 1777 8823
rect 1636 8792 1777 8820
rect 1636 8780 1642 8792
rect 1765 8789 1777 8792
rect 1811 8789 1823 8823
rect 1765 8783 1823 8789
rect 1854 8780 1860 8832
rect 1912 8820 1918 8832
rect 2682 8820 2688 8832
rect 1912 8792 2688 8820
rect 1912 8780 1918 8792
rect 2682 8780 2688 8792
rect 2740 8780 2746 8832
rect 2774 8780 2780 8832
rect 2832 8820 2838 8832
rect 4154 8820 4160 8832
rect 2832 8792 4160 8820
rect 2832 8780 2838 8792
rect 4154 8780 4160 8792
rect 4212 8780 4218 8832
rect 4246 8780 4252 8832
rect 4304 8780 4310 8832
rect 4890 8780 4896 8832
rect 4948 8780 4954 8832
rect 5350 8780 5356 8832
rect 5408 8780 5414 8832
rect 7190 8780 7196 8832
rect 7248 8820 7254 8832
rect 7834 8820 7840 8832
rect 7248 8792 7840 8820
rect 7248 8780 7254 8792
rect 7834 8780 7840 8792
rect 7892 8780 7898 8832
rect 8202 8780 8208 8832
rect 8260 8820 8266 8832
rect 10060 8820 10088 8996
rect 10318 8984 10324 8996
rect 10376 8984 10382 9036
rect 11606 8984 11612 9036
rect 11664 9024 11670 9036
rect 12618 9024 12624 9036
rect 11664 8996 12624 9024
rect 11664 8984 11670 8996
rect 12618 8984 12624 8996
rect 12676 9024 12682 9036
rect 16316 9024 16344 9064
rect 16758 9052 16764 9064
rect 16816 9092 16822 9104
rect 16816 9064 16991 9092
rect 16816 9052 16822 9064
rect 12676 8996 16344 9024
rect 12676 8984 12682 8996
rect 16390 8984 16396 9036
rect 16448 9024 16454 9036
rect 16485 9027 16543 9033
rect 16485 9024 16497 9027
rect 16448 8996 16497 9024
rect 16448 8984 16454 8996
rect 16485 8993 16497 8996
rect 16531 8993 16543 9027
rect 16485 8987 16543 8993
rect 16963 9024 16991 9064
rect 17218 9052 17224 9104
rect 17276 9092 17282 9104
rect 18690 9092 18696 9104
rect 17276 9064 18696 9092
rect 17276 9052 17282 9064
rect 18690 9052 18696 9064
rect 18748 9052 18754 9104
rect 16963 8996 17724 9024
rect 10134 8916 10140 8968
rect 10192 8956 10198 8968
rect 10192 8928 11192 8956
rect 10192 8916 10198 8928
rect 10318 8848 10324 8900
rect 10376 8888 10382 8900
rect 11164 8897 11192 8928
rect 12802 8916 12808 8968
rect 12860 8956 12866 8968
rect 13630 8956 13636 8968
rect 12860 8928 13636 8956
rect 12860 8916 12866 8928
rect 13630 8916 13636 8928
rect 13688 8916 13694 8968
rect 13998 8916 14004 8968
rect 14056 8956 14062 8968
rect 14182 8956 14188 8968
rect 14056 8928 14188 8956
rect 14056 8916 14062 8928
rect 14182 8916 14188 8928
rect 14240 8916 14246 8968
rect 16577 8959 16635 8965
rect 16577 8925 16589 8959
rect 16623 8956 16635 8959
rect 16666 8956 16672 8968
rect 16623 8928 16672 8956
rect 16623 8925 16635 8928
rect 16577 8919 16635 8925
rect 16666 8916 16672 8928
rect 16724 8916 16730 8968
rect 16963 8965 16991 8996
rect 16948 8959 17006 8965
rect 16948 8925 16960 8959
rect 16994 8925 17006 8959
rect 17218 8956 17224 8968
rect 16948 8919 17006 8925
rect 17052 8928 17224 8956
rect 10933 8891 10991 8897
rect 10933 8888 10945 8891
rect 10376 8860 10945 8888
rect 10376 8848 10382 8860
rect 10933 8857 10945 8860
rect 10979 8857 10991 8891
rect 10933 8851 10991 8857
rect 11149 8891 11207 8897
rect 11149 8857 11161 8891
rect 11195 8857 11207 8891
rect 11149 8851 11207 8857
rect 12526 8848 12532 8900
rect 12584 8888 12590 8900
rect 16482 8888 16488 8900
rect 12584 8860 16488 8888
rect 12584 8848 12590 8860
rect 16482 8848 16488 8860
rect 16540 8848 16546 8900
rect 17052 8888 17080 8928
rect 17218 8916 17224 8928
rect 17276 8956 17282 8968
rect 17696 8965 17724 8996
rect 17497 8959 17555 8965
rect 17497 8956 17509 8959
rect 17276 8928 17509 8956
rect 17276 8916 17282 8928
rect 17497 8925 17509 8928
rect 17543 8925 17555 8959
rect 17497 8919 17555 8925
rect 17681 8959 17739 8965
rect 17681 8925 17693 8959
rect 17727 8925 17739 8959
rect 17681 8919 17739 8925
rect 18233 8959 18291 8965
rect 18233 8925 18245 8959
rect 18279 8925 18291 8959
rect 18233 8919 18291 8925
rect 18248 8888 18276 8919
rect 16700 8860 17080 8888
rect 17144 8860 18276 8888
rect 8260 8792 10088 8820
rect 8260 8780 8266 8792
rect 10410 8780 10416 8832
rect 10468 8780 10474 8832
rect 11882 8780 11888 8832
rect 11940 8820 11946 8832
rect 12894 8820 12900 8832
rect 11940 8792 12900 8820
rect 11940 8780 11946 8792
rect 12894 8780 12900 8792
rect 12952 8820 12958 8832
rect 15102 8820 15108 8832
rect 12952 8792 15108 8820
rect 12952 8780 12958 8792
rect 15102 8780 15108 8792
rect 15160 8780 15166 8832
rect 16390 8780 16396 8832
rect 16448 8820 16454 8832
rect 16700 8820 16728 8860
rect 16448 8792 16728 8820
rect 16448 8780 16454 8792
rect 16758 8780 16764 8832
rect 16816 8820 16822 8832
rect 17144 8829 17172 8860
rect 16945 8823 17003 8829
rect 16945 8820 16957 8823
rect 16816 8792 16957 8820
rect 16816 8780 16822 8792
rect 16945 8789 16957 8792
rect 16991 8789 17003 8823
rect 16945 8783 17003 8789
rect 17129 8823 17187 8829
rect 17129 8789 17141 8823
rect 17175 8789 17187 8823
rect 17129 8783 17187 8789
rect 17589 8823 17647 8829
rect 17589 8789 17601 8823
rect 17635 8820 17647 8823
rect 17954 8820 17960 8832
rect 17635 8792 17960 8820
rect 17635 8789 17647 8792
rect 17589 8783 17647 8789
rect 17954 8780 17960 8792
rect 18012 8780 18018 8832
rect 18414 8780 18420 8832
rect 18472 8780 18478 8832
rect 1104 8730 18860 8752
rect 1104 8678 2610 8730
rect 2662 8678 2674 8730
rect 2726 8678 2738 8730
rect 2790 8678 2802 8730
rect 2854 8678 2866 8730
rect 2918 8678 7610 8730
rect 7662 8678 7674 8730
rect 7726 8678 7738 8730
rect 7790 8678 7802 8730
rect 7854 8678 7866 8730
rect 7918 8678 12610 8730
rect 12662 8678 12674 8730
rect 12726 8678 12738 8730
rect 12790 8678 12802 8730
rect 12854 8678 12866 8730
rect 12918 8678 17610 8730
rect 17662 8678 17674 8730
rect 17726 8678 17738 8730
rect 17790 8678 17802 8730
rect 17854 8678 17866 8730
rect 17918 8678 18860 8730
rect 1104 8656 18860 8678
rect 1118 8576 1124 8628
rect 1176 8616 1182 8628
rect 1670 8616 1676 8628
rect 1176 8588 1676 8616
rect 1176 8576 1182 8588
rect 1670 8576 1676 8588
rect 1728 8576 1734 8628
rect 2130 8576 2136 8628
rect 2188 8576 2194 8628
rect 2222 8576 2228 8628
rect 2280 8616 2286 8628
rect 2317 8619 2375 8625
rect 2317 8616 2329 8619
rect 2280 8588 2329 8616
rect 2280 8576 2286 8588
rect 2317 8585 2329 8588
rect 2363 8585 2375 8619
rect 2317 8579 2375 8585
rect 2406 8576 2412 8628
rect 2464 8616 2470 8628
rect 2590 8616 2596 8628
rect 2464 8588 2596 8616
rect 2464 8576 2470 8588
rect 2590 8576 2596 8588
rect 2648 8576 2654 8628
rect 3878 8616 3884 8628
rect 2746 8588 3884 8616
rect 1762 8508 1768 8560
rect 1820 8548 1826 8560
rect 1949 8551 2007 8557
rect 1949 8548 1961 8551
rect 1820 8520 1961 8548
rect 1820 8508 1826 8520
rect 1949 8517 1961 8520
rect 1995 8517 2007 8551
rect 2746 8548 2774 8588
rect 3878 8576 3884 8588
rect 3936 8576 3942 8628
rect 4246 8576 4252 8628
rect 4304 8616 4310 8628
rect 5258 8616 5264 8628
rect 4304 8588 5264 8616
rect 4304 8576 4310 8588
rect 5258 8576 5264 8588
rect 5316 8576 5322 8628
rect 5994 8576 6000 8628
rect 6052 8616 6058 8628
rect 7009 8619 7067 8625
rect 7009 8616 7021 8619
rect 6052 8588 7021 8616
rect 6052 8576 6058 8588
rect 7009 8585 7021 8588
rect 7055 8585 7067 8619
rect 7009 8579 7067 8585
rect 7098 8576 7104 8628
rect 7156 8616 7162 8628
rect 7650 8616 7656 8628
rect 7156 8588 7656 8616
rect 7156 8576 7162 8588
rect 7650 8576 7656 8588
rect 7708 8576 7714 8628
rect 7742 8576 7748 8628
rect 7800 8616 7806 8628
rect 8662 8616 8668 8628
rect 7800 8588 8668 8616
rect 7800 8576 7806 8588
rect 8662 8576 8668 8588
rect 8720 8616 8726 8628
rect 9401 8619 9459 8625
rect 9401 8616 9413 8619
rect 8720 8588 9413 8616
rect 8720 8576 8726 8588
rect 9401 8585 9413 8588
rect 9447 8585 9459 8619
rect 10045 8619 10103 8625
rect 9401 8579 9459 8585
rect 9508 8588 9996 8616
rect 3418 8548 3424 8560
rect 1949 8511 2007 8517
rect 2148 8520 2774 8548
rect 3068 8520 3424 8548
rect 1670 8440 1676 8492
rect 1728 8480 1734 8492
rect 2148 8480 2176 8520
rect 1728 8452 2176 8480
rect 2225 8483 2283 8489
rect 1728 8440 1734 8452
rect 2225 8449 2237 8483
rect 2271 8449 2283 8483
rect 2225 8443 2283 8449
rect 198 8372 204 8424
rect 256 8412 262 8424
rect 2240 8412 2268 8443
rect 2406 8440 2412 8492
rect 2464 8480 2470 8492
rect 3068 8489 3096 8520
rect 3418 8508 3424 8520
rect 3476 8508 3482 8560
rect 4525 8551 4583 8557
rect 3620 8520 4200 8548
rect 3053 8483 3111 8489
rect 3053 8480 3065 8483
rect 2464 8452 3065 8480
rect 2464 8440 2470 8452
rect 3053 8449 3065 8452
rect 3099 8449 3111 8483
rect 3053 8443 3111 8449
rect 3145 8483 3203 8489
rect 3145 8449 3157 8483
rect 3191 8449 3203 8483
rect 3145 8443 3203 8449
rect 2314 8412 2320 8424
rect 256 8384 2320 8412
rect 256 8372 262 8384
rect 2314 8372 2320 8384
rect 2372 8372 2378 8424
rect 2590 8372 2596 8424
rect 2648 8372 2654 8424
rect 2958 8372 2964 8424
rect 3016 8412 3022 8424
rect 3160 8412 3188 8443
rect 3510 8440 3516 8492
rect 3568 8480 3574 8492
rect 3620 8480 3648 8520
rect 3568 8466 3648 8480
rect 3568 8452 3634 8466
rect 3568 8440 3574 8452
rect 3016 8384 3188 8412
rect 3734 8415 3792 8421
rect 3016 8372 3022 8384
rect 3734 8381 3746 8415
rect 3780 8412 3792 8415
rect 3878 8412 3884 8424
rect 3780 8384 3884 8412
rect 3780 8381 3792 8384
rect 3734 8375 3792 8381
rect 3878 8372 3884 8384
rect 3936 8372 3942 8424
rect 4172 8412 4200 8520
rect 4525 8517 4537 8551
rect 4571 8548 4583 8551
rect 4706 8548 4712 8560
rect 4571 8520 4712 8548
rect 4571 8517 4583 8520
rect 4525 8511 4583 8517
rect 4706 8508 4712 8520
rect 4764 8508 4770 8560
rect 9508 8548 9536 8588
rect 5000 8520 9536 8548
rect 4246 8440 4252 8492
rect 4304 8480 4310 8492
rect 5000 8489 5028 8520
rect 4801 8483 4859 8489
rect 4801 8480 4813 8483
rect 4304 8452 4813 8480
rect 4304 8440 4310 8452
rect 4801 8449 4813 8452
rect 4847 8449 4859 8483
rect 4801 8443 4859 8449
rect 4985 8483 5043 8489
rect 4985 8449 4997 8483
rect 5031 8449 5043 8483
rect 4985 8443 5043 8449
rect 5353 8483 5411 8489
rect 5353 8449 5365 8483
rect 5399 8449 5411 8483
rect 5353 8443 5411 8449
rect 5537 8483 5595 8489
rect 5537 8449 5549 8483
rect 5583 8480 5595 8483
rect 5718 8480 5724 8492
rect 5583 8452 5724 8480
rect 5583 8449 5595 8452
rect 5537 8443 5595 8449
rect 5258 8412 5264 8424
rect 4172 8384 5264 8412
rect 5258 8372 5264 8384
rect 5316 8412 5322 8424
rect 5368 8412 5396 8443
rect 5718 8440 5724 8452
rect 5776 8440 5782 8492
rect 6365 8483 6423 8489
rect 6365 8449 6377 8483
rect 6411 8480 6423 8483
rect 6454 8480 6460 8492
rect 6411 8452 6460 8480
rect 6411 8449 6423 8452
rect 6365 8443 6423 8449
rect 6454 8440 6460 8452
rect 6512 8440 6518 8492
rect 6546 8440 6552 8492
rect 6604 8440 6610 8492
rect 6641 8483 6699 8489
rect 6641 8449 6653 8483
rect 6687 8449 6699 8483
rect 6641 8443 6699 8449
rect 5316 8384 5396 8412
rect 5316 8372 5322 8384
rect 5994 8372 6000 8424
rect 6052 8372 6058 8424
rect 2222 8304 2228 8356
rect 2280 8344 2286 8356
rect 2501 8347 2559 8353
rect 2280 8316 2452 8344
rect 2280 8304 2286 8316
rect 2038 8236 2044 8288
rect 2096 8276 2102 8288
rect 2314 8276 2320 8288
rect 2096 8248 2320 8276
rect 2096 8236 2102 8248
rect 2314 8236 2320 8248
rect 2372 8236 2378 8288
rect 2424 8276 2452 8316
rect 2501 8313 2513 8347
rect 2547 8344 2559 8347
rect 4338 8344 4344 8356
rect 2547 8316 4344 8344
rect 2547 8313 2559 8316
rect 2501 8307 2559 8313
rect 4338 8304 4344 8316
rect 4396 8304 4402 8356
rect 4798 8304 4804 8356
rect 4856 8344 4862 8356
rect 6656 8344 6684 8443
rect 6730 8440 6736 8492
rect 6788 8440 6794 8492
rect 6822 8440 6828 8492
rect 6880 8480 6886 8492
rect 7193 8483 7251 8489
rect 7193 8480 7205 8483
rect 6880 8452 7205 8480
rect 6880 8440 6886 8452
rect 7193 8449 7205 8452
rect 7239 8449 7251 8483
rect 7193 8443 7251 8449
rect 7377 8483 7435 8489
rect 7377 8449 7389 8483
rect 7423 8480 7435 8483
rect 7558 8480 7564 8492
rect 7423 8452 7564 8480
rect 7423 8449 7435 8452
rect 7377 8443 7435 8449
rect 7558 8440 7564 8452
rect 7616 8440 7622 8492
rect 7650 8440 7656 8492
rect 7708 8480 7714 8492
rect 8570 8480 8576 8492
rect 7708 8452 8576 8480
rect 7708 8440 7714 8452
rect 8570 8440 8576 8452
rect 8628 8440 8634 8492
rect 8662 8440 8668 8492
rect 8720 8480 8726 8492
rect 9306 8480 9312 8492
rect 8720 8452 9312 8480
rect 8720 8440 8726 8452
rect 9306 8440 9312 8452
rect 9364 8440 9370 8492
rect 9582 8440 9588 8492
rect 9640 8480 9646 8492
rect 9968 8480 9996 8588
rect 10045 8585 10057 8619
rect 10091 8585 10103 8619
rect 10045 8579 10103 8585
rect 10060 8548 10088 8579
rect 10134 8576 10140 8628
rect 10192 8616 10198 8628
rect 10413 8619 10471 8625
rect 10413 8616 10425 8619
rect 10192 8588 10425 8616
rect 10192 8576 10198 8588
rect 10413 8585 10425 8588
rect 10459 8585 10471 8619
rect 10413 8579 10471 8585
rect 10686 8576 10692 8628
rect 10744 8616 10750 8628
rect 13170 8616 13176 8628
rect 10744 8588 13176 8616
rect 10744 8576 10750 8588
rect 13170 8576 13176 8588
rect 13228 8576 13234 8628
rect 15102 8576 15108 8628
rect 15160 8616 15166 8628
rect 16390 8616 16396 8628
rect 15160 8588 16396 8616
rect 15160 8576 15166 8588
rect 16390 8576 16396 8588
rect 16448 8576 16454 8628
rect 10597 8551 10655 8557
rect 10060 8520 10548 8548
rect 10137 8483 10195 8489
rect 10137 8480 10149 8483
rect 9640 8452 9904 8480
rect 9968 8452 10149 8480
rect 9640 8440 9646 8452
rect 6748 8412 6776 8440
rect 7834 8412 7840 8424
rect 6748 8384 7840 8412
rect 7834 8372 7840 8384
rect 7892 8372 7898 8424
rect 9766 8412 9772 8424
rect 8266 8384 9772 8412
rect 4856 8316 6684 8344
rect 6917 8347 6975 8353
rect 4856 8304 4862 8316
rect 6917 8313 6929 8347
rect 6963 8344 6975 8347
rect 8266 8344 8294 8384
rect 9766 8372 9772 8384
rect 9824 8372 9830 8424
rect 6963 8316 8294 8344
rect 6963 8313 6975 8316
rect 6917 8307 6975 8313
rect 8570 8304 8576 8356
rect 8628 8344 8634 8356
rect 9876 8344 9904 8452
rect 10137 8449 10149 8452
rect 10183 8449 10195 8483
rect 10137 8443 10195 8449
rect 8628 8316 9904 8344
rect 10152 8344 10180 8443
rect 10318 8440 10324 8492
rect 10376 8440 10382 8492
rect 10520 8480 10548 8520
rect 10597 8517 10609 8551
rect 10643 8548 10655 8551
rect 11330 8548 11336 8560
rect 10643 8520 11336 8548
rect 10643 8517 10655 8520
rect 10597 8511 10655 8517
rect 11330 8508 11336 8520
rect 11388 8508 11394 8560
rect 12158 8508 12164 8560
rect 12216 8548 12222 8560
rect 13722 8548 13728 8560
rect 12216 8520 13728 8548
rect 12216 8508 12222 8520
rect 13722 8508 13728 8520
rect 13780 8508 13786 8560
rect 13998 8508 14004 8560
rect 14056 8548 14062 8560
rect 15746 8548 15752 8560
rect 14056 8520 15752 8548
rect 14056 8508 14062 8520
rect 15746 8508 15752 8520
rect 15804 8508 15810 8560
rect 18782 8548 18788 8560
rect 16960 8520 18788 8548
rect 10962 8480 10968 8492
rect 10520 8452 10968 8480
rect 10962 8440 10968 8452
rect 11020 8440 11026 8492
rect 12250 8440 12256 8492
rect 12308 8480 12314 8492
rect 15378 8480 15384 8492
rect 12308 8452 15384 8480
rect 12308 8440 12314 8452
rect 15378 8440 15384 8452
rect 15436 8480 15442 8492
rect 16960 8489 16988 8520
rect 18782 8508 18788 8520
rect 18840 8508 18846 8560
rect 16669 8483 16727 8489
rect 16669 8480 16681 8483
rect 15436 8452 16681 8480
rect 15436 8440 15442 8452
rect 16669 8449 16681 8452
rect 16715 8449 16727 8483
rect 16669 8443 16727 8449
rect 16945 8483 17003 8489
rect 16945 8449 16957 8483
rect 16991 8449 17003 8483
rect 16945 8443 17003 8449
rect 17037 8483 17095 8489
rect 17037 8449 17049 8483
rect 17083 8480 17095 8483
rect 18046 8480 18052 8492
rect 17083 8452 18052 8480
rect 17083 8449 17095 8452
rect 17037 8443 17095 8449
rect 18046 8440 18052 8452
rect 18104 8440 18110 8492
rect 10226 8372 10232 8424
rect 10284 8412 10290 8424
rect 15470 8412 15476 8424
rect 10284 8384 15476 8412
rect 10284 8372 10290 8384
rect 15470 8372 15476 8384
rect 15528 8372 15534 8424
rect 15654 8372 15660 8424
rect 15712 8412 15718 8424
rect 19518 8412 19524 8424
rect 15712 8384 19524 8412
rect 15712 8372 15718 8384
rect 19518 8372 19524 8384
rect 19576 8372 19582 8424
rect 10410 8344 10416 8356
rect 10152 8316 10416 8344
rect 8628 8304 8634 8316
rect 10410 8304 10416 8316
rect 10468 8304 10474 8356
rect 10594 8304 10600 8356
rect 10652 8304 10658 8356
rect 11330 8304 11336 8356
rect 11388 8344 11394 8356
rect 11388 8316 12940 8344
rect 11388 8304 11394 8316
rect 2682 8276 2688 8288
rect 2424 8248 2688 8276
rect 2682 8236 2688 8248
rect 2740 8236 2746 8288
rect 3050 8236 3056 8288
rect 3108 8276 3114 8288
rect 3329 8279 3387 8285
rect 3329 8276 3341 8279
rect 3108 8248 3341 8276
rect 3108 8236 3114 8248
rect 3329 8245 3341 8248
rect 3375 8245 3387 8279
rect 3329 8239 3387 8245
rect 5074 8236 5080 8288
rect 5132 8276 5138 8288
rect 5534 8276 5540 8288
rect 5132 8248 5540 8276
rect 5132 8236 5138 8248
rect 5534 8236 5540 8248
rect 5592 8236 5598 8288
rect 7006 8236 7012 8288
rect 7064 8276 7070 8288
rect 8110 8276 8116 8288
rect 7064 8248 8116 8276
rect 7064 8236 7070 8248
rect 8110 8236 8116 8248
rect 8168 8236 8174 8288
rect 8754 8236 8760 8288
rect 8812 8276 8818 8288
rect 9306 8276 9312 8288
rect 8812 8248 9312 8276
rect 8812 8236 8818 8248
rect 9306 8236 9312 8248
rect 9364 8236 9370 8288
rect 9398 8236 9404 8288
rect 9456 8276 9462 8288
rect 9674 8276 9680 8288
rect 9456 8248 9680 8276
rect 9456 8236 9462 8248
rect 9674 8236 9680 8248
rect 9732 8236 9738 8288
rect 9950 8236 9956 8288
rect 10008 8276 10014 8288
rect 10686 8276 10692 8288
rect 10008 8248 10692 8276
rect 10008 8236 10014 8248
rect 10686 8236 10692 8248
rect 10744 8236 10750 8288
rect 11146 8236 11152 8288
rect 11204 8276 11210 8288
rect 12802 8276 12808 8288
rect 11204 8248 12808 8276
rect 11204 8236 11210 8248
rect 12802 8236 12808 8248
rect 12860 8236 12866 8288
rect 12912 8276 12940 8316
rect 13722 8304 13728 8356
rect 13780 8344 13786 8356
rect 14550 8344 14556 8356
rect 13780 8316 14556 8344
rect 13780 8304 13786 8316
rect 14550 8304 14556 8316
rect 14608 8304 14614 8356
rect 14918 8276 14924 8288
rect 12912 8248 14924 8276
rect 14918 8236 14924 8248
rect 14976 8236 14982 8288
rect 15470 8236 15476 8288
rect 15528 8276 15534 8288
rect 16761 8279 16819 8285
rect 16761 8276 16773 8279
rect 15528 8248 16773 8276
rect 15528 8236 15534 8248
rect 16761 8245 16773 8248
rect 16807 8245 16819 8279
rect 16761 8239 16819 8245
rect 17221 8279 17279 8285
rect 17221 8245 17233 8279
rect 17267 8276 17279 8279
rect 17586 8276 17592 8288
rect 17267 8248 17592 8276
rect 17267 8245 17279 8248
rect 17221 8239 17279 8245
rect 17586 8236 17592 8248
rect 17644 8236 17650 8288
rect 1104 8186 18860 8208
rect 1104 8134 1950 8186
rect 2002 8134 2014 8186
rect 2066 8134 2078 8186
rect 2130 8134 2142 8186
rect 2194 8134 2206 8186
rect 2258 8134 6950 8186
rect 7002 8134 7014 8186
rect 7066 8134 7078 8186
rect 7130 8134 7142 8186
rect 7194 8134 7206 8186
rect 7258 8134 11950 8186
rect 12002 8134 12014 8186
rect 12066 8134 12078 8186
rect 12130 8134 12142 8186
rect 12194 8134 12206 8186
rect 12258 8134 16950 8186
rect 17002 8134 17014 8186
rect 17066 8134 17078 8186
rect 17130 8134 17142 8186
rect 17194 8134 17206 8186
rect 17258 8134 18860 8186
rect 1104 8112 18860 8134
rect 2774 8032 2780 8084
rect 2832 8072 2838 8084
rect 4614 8072 4620 8084
rect 2832 8044 4620 8072
rect 2832 8032 2838 8044
rect 4614 8032 4620 8044
rect 4672 8032 4678 8084
rect 5258 8032 5264 8084
rect 5316 8072 5322 8084
rect 5997 8075 6055 8081
rect 5997 8072 6009 8075
rect 5316 8044 6009 8072
rect 5316 8032 5322 8044
rect 5997 8041 6009 8044
rect 6043 8041 6055 8075
rect 12434 8072 12440 8084
rect 5997 8035 6055 8041
rect 6372 8044 12440 8072
rect 750 7964 756 8016
rect 808 8004 814 8016
rect 1673 8007 1731 8013
rect 1673 8004 1685 8007
rect 808 7976 1685 8004
rect 808 7964 814 7976
rect 1673 7973 1685 7976
rect 1719 7973 1731 8007
rect 1673 7967 1731 7973
rect 2501 8007 2559 8013
rect 2501 7973 2513 8007
rect 2547 8004 2559 8007
rect 2866 8004 2872 8016
rect 2547 7976 2872 8004
rect 2547 7973 2559 7976
rect 2501 7967 2559 7973
rect 1688 7936 1716 7967
rect 2866 7964 2872 7976
rect 2924 7964 2930 8016
rect 6270 8004 6276 8016
rect 3528 7976 6276 8004
rect 3528 7936 3556 7976
rect 6270 7964 6276 7976
rect 6328 7964 6334 8016
rect 1688 7908 3556 7936
rect 3602 7896 3608 7948
rect 3660 7936 3666 7948
rect 3878 7936 3884 7948
rect 3660 7908 3884 7936
rect 3660 7896 3666 7908
rect 3878 7896 3884 7908
rect 3936 7936 3942 7948
rect 6372 7936 6400 8044
rect 12434 8032 12440 8044
rect 12492 8032 12498 8084
rect 13103 8075 13161 8081
rect 13103 8041 13115 8075
rect 13149 8072 13161 8075
rect 13906 8072 13912 8084
rect 13149 8044 13912 8072
rect 13149 8041 13161 8044
rect 13103 8035 13161 8041
rect 13906 8032 13912 8044
rect 13964 8032 13970 8084
rect 15749 8075 15807 8081
rect 15749 8041 15761 8075
rect 15795 8072 15807 8075
rect 16022 8072 16028 8084
rect 15795 8044 16028 8072
rect 15795 8041 15807 8044
rect 15749 8035 15807 8041
rect 16022 8032 16028 8044
rect 16080 8032 16086 8084
rect 16758 8072 16764 8084
rect 16132 8044 16764 8072
rect 11238 8004 11244 8016
rect 3936 7908 6400 7936
rect 6472 7976 8064 8004
rect 3936 7896 3942 7908
rect 1397 7871 1455 7877
rect 1397 7837 1409 7871
rect 1443 7868 1455 7871
rect 1443 7840 4479 7868
rect 1443 7837 1455 7840
rect 1397 7831 1455 7837
rect 1762 7760 1768 7812
rect 1820 7800 1826 7812
rect 2685 7803 2743 7809
rect 2685 7800 2697 7803
rect 1820 7772 2697 7800
rect 1820 7760 1826 7772
rect 2685 7769 2697 7772
rect 2731 7769 2743 7803
rect 2685 7763 2743 7769
rect 2869 7803 2927 7809
rect 2869 7769 2881 7803
rect 2915 7800 2927 7803
rect 3878 7800 3884 7812
rect 2915 7772 3884 7800
rect 2915 7769 2927 7772
rect 2869 7763 2927 7769
rect 3878 7760 3884 7772
rect 3936 7760 3942 7812
rect 4338 7760 4344 7812
rect 4396 7760 4402 7812
rect 1302 7692 1308 7744
rect 1360 7732 1366 7744
rect 1857 7735 1915 7741
rect 1857 7732 1869 7735
rect 1360 7704 1869 7732
rect 1360 7692 1366 7704
rect 1857 7701 1869 7704
rect 1903 7701 1915 7735
rect 1857 7695 1915 7701
rect 2774 7692 2780 7744
rect 2832 7732 2838 7744
rect 3050 7732 3056 7744
rect 2832 7704 3056 7732
rect 2832 7692 2838 7704
rect 3050 7692 3056 7704
rect 3108 7692 3114 7744
rect 4451 7732 4479 7840
rect 4522 7828 4528 7880
rect 4580 7828 4586 7880
rect 5828 7877 5856 7908
rect 5813 7871 5871 7877
rect 5813 7837 5825 7871
rect 5859 7837 5871 7871
rect 5813 7831 5871 7837
rect 5994 7828 6000 7880
rect 6052 7868 6058 7880
rect 6472 7868 6500 7976
rect 6638 7896 6644 7948
rect 6696 7936 6702 7948
rect 6696 7908 6868 7936
rect 6696 7896 6702 7908
rect 6052 7840 6500 7868
rect 6549 7871 6607 7877
rect 6052 7828 6058 7840
rect 6549 7837 6561 7871
rect 6595 7837 6607 7871
rect 6549 7831 6607 7837
rect 6564 7800 6592 7831
rect 6730 7828 6736 7880
rect 6788 7828 6794 7880
rect 6840 7877 6868 7908
rect 7190 7896 7196 7948
rect 7248 7896 7254 7948
rect 7282 7896 7288 7948
rect 7340 7936 7346 7948
rect 7926 7936 7932 7948
rect 7340 7908 7932 7936
rect 7340 7896 7346 7908
rect 7926 7896 7932 7908
rect 7984 7896 7990 7948
rect 8036 7936 8064 7976
rect 9416 7976 11244 8004
rect 9416 7936 9444 7976
rect 11238 7964 11244 7976
rect 11296 7964 11302 8016
rect 13265 8007 13323 8013
rect 13265 7973 13277 8007
rect 13311 8004 13323 8007
rect 13354 8004 13360 8016
rect 13311 7976 13360 8004
rect 13311 7973 13323 7976
rect 13265 7967 13323 7973
rect 13354 7964 13360 7976
rect 13412 7964 13418 8016
rect 15102 7964 15108 8016
rect 15160 8004 15166 8016
rect 15160 7976 15608 8004
rect 15160 7964 15166 7976
rect 8036 7908 9444 7936
rect 9677 7939 9735 7945
rect 9677 7905 9689 7939
rect 9723 7936 9735 7939
rect 9950 7936 9956 7948
rect 9723 7908 9956 7936
rect 9723 7905 9735 7908
rect 9677 7899 9735 7905
rect 9950 7896 9956 7908
rect 10008 7896 10014 7948
rect 10686 7896 10692 7948
rect 10744 7936 10750 7948
rect 12986 7936 12992 7948
rect 10744 7908 12992 7936
rect 10744 7896 10750 7908
rect 12986 7896 12992 7908
rect 13044 7896 13050 7948
rect 14476 7908 15332 7936
rect 6825 7871 6883 7877
rect 6825 7837 6837 7871
rect 6871 7837 6883 7871
rect 6825 7831 6883 7837
rect 6917 7871 6975 7877
rect 6917 7837 6929 7871
rect 6963 7868 6975 7871
rect 7558 7868 7564 7880
rect 6963 7840 7564 7868
rect 6963 7837 6975 7840
rect 6917 7831 6975 7837
rect 7558 7828 7564 7840
rect 7616 7828 7622 7880
rect 7834 7828 7840 7880
rect 7892 7868 7898 7880
rect 8202 7868 8208 7880
rect 7892 7840 8208 7868
rect 7892 7828 7898 7840
rect 8202 7828 8208 7840
rect 8260 7828 8266 7880
rect 8386 7828 8392 7880
rect 8444 7868 8450 7880
rect 8444 7840 9076 7868
rect 8444 7828 8450 7840
rect 6564 7772 7144 7800
rect 7006 7732 7012 7744
rect 4451 7704 7012 7732
rect 7006 7692 7012 7704
rect 7064 7692 7070 7744
rect 7116 7732 7144 7772
rect 7190 7760 7196 7812
rect 7248 7800 7254 7812
rect 9048 7800 9076 7840
rect 9122 7828 9128 7880
rect 9180 7868 9186 7880
rect 9217 7871 9275 7877
rect 9217 7868 9229 7871
rect 9180 7840 9229 7868
rect 9180 7828 9186 7840
rect 9217 7837 9229 7840
rect 9263 7837 9275 7871
rect 9217 7831 9275 7837
rect 9306 7828 9312 7880
rect 9364 7828 9370 7880
rect 9585 7871 9643 7877
rect 9585 7868 9597 7871
rect 9416 7840 9597 7868
rect 9416 7800 9444 7840
rect 9585 7837 9597 7840
rect 9631 7837 9643 7871
rect 9585 7831 9643 7837
rect 9766 7828 9772 7880
rect 9824 7828 9830 7880
rect 10778 7828 10784 7880
rect 10836 7828 10842 7880
rect 13814 7868 13820 7880
rect 12912 7840 13820 7868
rect 7248 7772 8984 7800
rect 9048 7772 9444 7800
rect 9493 7803 9551 7809
rect 7248 7760 7254 7772
rect 8110 7732 8116 7744
rect 7116 7704 8116 7732
rect 8110 7692 8116 7704
rect 8168 7692 8174 7744
rect 8956 7732 8984 7772
rect 9493 7769 9505 7803
rect 9539 7800 9551 7803
rect 10796 7800 10824 7828
rect 12912 7809 12940 7840
rect 13814 7828 13820 7840
rect 13872 7828 13878 7880
rect 13906 7828 13912 7880
rect 13964 7868 13970 7880
rect 14476 7868 14504 7908
rect 13964 7840 14504 7868
rect 13964 7828 13970 7840
rect 14826 7828 14832 7880
rect 14884 7868 14890 7880
rect 15105 7871 15163 7877
rect 15105 7868 15117 7871
rect 14884 7840 15117 7868
rect 14884 7828 14890 7840
rect 15105 7837 15117 7840
rect 15151 7837 15163 7871
rect 15105 7831 15163 7837
rect 15197 7871 15255 7877
rect 15197 7837 15209 7871
rect 15243 7837 15255 7871
rect 15197 7831 15255 7837
rect 9539 7772 10824 7800
rect 12897 7803 12955 7809
rect 9539 7769 9551 7772
rect 9493 7763 9551 7769
rect 12897 7769 12909 7803
rect 12943 7769 12955 7803
rect 12897 7763 12955 7769
rect 13113 7803 13171 7809
rect 13113 7769 13125 7803
rect 13159 7800 13171 7803
rect 13722 7800 13728 7812
rect 13159 7772 13728 7800
rect 13159 7769 13171 7772
rect 13113 7763 13171 7769
rect 13722 7760 13728 7772
rect 13780 7760 13786 7812
rect 10778 7732 10784 7744
rect 8956 7704 10784 7732
rect 10778 7692 10784 7704
rect 10836 7692 10842 7744
rect 11146 7692 11152 7744
rect 11204 7732 11210 7744
rect 11514 7732 11520 7744
rect 11204 7704 11520 7732
rect 11204 7692 11210 7704
rect 11514 7692 11520 7704
rect 11572 7732 11578 7744
rect 12618 7732 12624 7744
rect 11572 7704 12624 7732
rect 11572 7692 11578 7704
rect 12618 7692 12624 7704
rect 12676 7692 12682 7744
rect 12802 7692 12808 7744
rect 12860 7732 12866 7744
rect 13354 7732 13360 7744
rect 12860 7704 13360 7732
rect 12860 7692 12866 7704
rect 13354 7692 13360 7704
rect 13412 7692 13418 7744
rect 15212 7732 15240 7831
rect 15304 7800 15332 7908
rect 15378 7828 15384 7880
rect 15436 7828 15442 7880
rect 15470 7828 15476 7880
rect 15528 7828 15534 7880
rect 15580 7877 15608 7976
rect 15838 7964 15844 8016
rect 15896 8004 15902 8016
rect 16132 8004 16160 8044
rect 16758 8032 16764 8044
rect 16816 8032 16822 8084
rect 15896 7976 16160 8004
rect 15896 7964 15902 7976
rect 16206 7936 16212 7948
rect 15948 7908 16212 7936
rect 15948 7877 15976 7908
rect 16206 7896 16212 7908
rect 16264 7896 16270 7948
rect 15565 7871 15623 7877
rect 15565 7837 15577 7871
rect 15611 7837 15623 7871
rect 15565 7831 15623 7837
rect 15841 7871 15899 7877
rect 15841 7837 15853 7871
rect 15887 7837 15899 7871
rect 15841 7831 15899 7837
rect 15933 7871 15991 7877
rect 15933 7837 15945 7871
rect 15979 7837 15991 7871
rect 15933 7831 15991 7837
rect 15856 7800 15884 7831
rect 16114 7828 16120 7880
rect 16172 7828 16178 7880
rect 17034 7828 17040 7880
rect 17092 7868 17098 7880
rect 17497 7871 17555 7877
rect 17497 7868 17509 7871
rect 17092 7840 17509 7868
rect 17092 7828 17098 7840
rect 17497 7837 17509 7840
rect 17543 7837 17555 7871
rect 17497 7831 17555 7837
rect 18049 7871 18107 7877
rect 18049 7837 18061 7871
rect 18095 7868 18107 7871
rect 18138 7868 18144 7880
rect 18095 7840 18144 7868
rect 18095 7837 18107 7840
rect 18049 7831 18107 7837
rect 18138 7828 18144 7840
rect 18196 7828 18202 7880
rect 15304 7772 15884 7800
rect 17218 7760 17224 7812
rect 17276 7800 17282 7812
rect 17313 7803 17371 7809
rect 17313 7800 17325 7803
rect 17276 7772 17325 7800
rect 17276 7760 17282 7772
rect 17313 7769 17325 7772
rect 17359 7800 17371 7803
rect 19058 7800 19064 7812
rect 17359 7772 19064 7800
rect 17359 7769 17371 7772
rect 17313 7763 17371 7769
rect 19058 7760 19064 7772
rect 19116 7760 19122 7812
rect 15838 7732 15844 7744
rect 15212 7704 15844 7732
rect 15838 7692 15844 7704
rect 15896 7692 15902 7744
rect 16298 7692 16304 7744
rect 16356 7692 16362 7744
rect 1104 7642 18860 7664
rect 1104 7590 2610 7642
rect 2662 7590 2674 7642
rect 2726 7590 2738 7642
rect 2790 7590 2802 7642
rect 2854 7590 2866 7642
rect 2918 7590 7610 7642
rect 7662 7590 7674 7642
rect 7726 7590 7738 7642
rect 7790 7590 7802 7642
rect 7854 7590 7866 7642
rect 7918 7590 12610 7642
rect 12662 7590 12674 7642
rect 12726 7590 12738 7642
rect 12790 7590 12802 7642
rect 12854 7590 12866 7642
rect 12918 7590 17610 7642
rect 17662 7590 17674 7642
rect 17726 7590 17738 7642
rect 17790 7590 17802 7642
rect 17854 7590 17866 7642
rect 17918 7590 18860 7642
rect 1104 7568 18860 7590
rect 4706 7488 4712 7540
rect 4764 7528 4770 7540
rect 5258 7528 5264 7540
rect 4764 7500 5264 7528
rect 4764 7488 4770 7500
rect 5258 7488 5264 7500
rect 5316 7528 5322 7540
rect 8386 7528 8392 7540
rect 5316 7500 8392 7528
rect 5316 7488 5322 7500
rect 8386 7488 8392 7500
rect 8444 7488 8450 7540
rect 8846 7488 8852 7540
rect 8904 7528 8910 7540
rect 9401 7531 9459 7537
rect 9401 7528 9413 7531
rect 8904 7500 9413 7528
rect 8904 7488 8910 7500
rect 9401 7497 9413 7500
rect 9447 7497 9459 7531
rect 9401 7491 9459 7497
rect 9582 7488 9588 7540
rect 9640 7528 9646 7540
rect 9766 7528 9772 7540
rect 9640 7500 9772 7528
rect 9640 7488 9646 7500
rect 9766 7488 9772 7500
rect 9824 7528 9830 7540
rect 10594 7528 10600 7540
rect 9824 7500 10600 7528
rect 9824 7488 9830 7500
rect 10594 7488 10600 7500
rect 10652 7488 10658 7540
rect 10870 7488 10876 7540
rect 10928 7488 10934 7540
rect 11514 7488 11520 7540
rect 11572 7528 11578 7540
rect 13078 7528 13084 7540
rect 11572 7500 13084 7528
rect 11572 7488 11578 7500
rect 13078 7488 13084 7500
rect 13136 7488 13142 7540
rect 16298 7528 16304 7540
rect 14108 7500 16304 7528
rect 1486 7420 1492 7472
rect 1544 7460 1550 7472
rect 4890 7460 4896 7472
rect 1544 7432 4896 7460
rect 1544 7420 1550 7432
rect 4890 7420 4896 7432
rect 4948 7420 4954 7472
rect 6270 7420 6276 7472
rect 6328 7460 6334 7472
rect 8205 7463 8263 7469
rect 6328 7432 7788 7460
rect 6328 7420 6334 7432
rect 4338 7392 4344 7404
rect 4264 7364 4344 7392
rect 4264 7333 4292 7364
rect 4338 7352 4344 7364
rect 4396 7392 4402 7404
rect 7469 7398 7527 7401
rect 7392 7395 7527 7398
rect 7392 7392 7481 7395
rect 4396 7370 7481 7392
rect 4396 7364 7420 7370
rect 4396 7352 4402 7364
rect 7469 7361 7481 7370
rect 7515 7361 7527 7395
rect 7469 7355 7527 7361
rect 7558 7352 7564 7404
rect 7616 7352 7622 7404
rect 7760 7401 7788 7432
rect 8205 7429 8217 7463
rect 8251 7460 8263 7463
rect 8294 7460 8300 7472
rect 8251 7432 8300 7460
rect 8251 7429 8263 7432
rect 8205 7423 8263 7429
rect 8294 7420 8300 7432
rect 8352 7420 8358 7472
rect 10888 7460 10916 7488
rect 8772 7432 10916 7460
rect 7745 7395 7803 7401
rect 7745 7361 7757 7395
rect 7791 7361 7803 7395
rect 7745 7355 7803 7361
rect 4249 7327 4307 7333
rect 4249 7293 4261 7327
rect 4295 7293 4307 7327
rect 4249 7287 4307 7293
rect 4522 7284 4528 7336
rect 4580 7284 4586 7336
rect 6270 7284 6276 7336
rect 6328 7324 6334 7336
rect 6914 7324 6920 7336
rect 6328 7296 6920 7324
rect 6328 7284 6334 7296
rect 6914 7284 6920 7296
rect 6972 7284 6978 7336
rect 7098 7284 7104 7336
rect 7156 7324 7162 7336
rect 7650 7324 7656 7336
rect 7156 7296 7656 7324
rect 7156 7284 7162 7296
rect 7650 7284 7656 7296
rect 7708 7284 7714 7336
rect 7760 7324 7788 7355
rect 8110 7352 8116 7404
rect 8168 7392 8174 7404
rect 8662 7392 8668 7404
rect 8168 7364 8668 7392
rect 8168 7352 8174 7364
rect 8662 7352 8668 7364
rect 8720 7352 8726 7404
rect 8772 7401 8800 7432
rect 11054 7420 11060 7472
rect 11112 7460 11118 7472
rect 14108 7460 14136 7500
rect 16298 7488 16304 7500
rect 16356 7488 16362 7540
rect 11112 7432 14136 7460
rect 11112 7420 11118 7432
rect 15102 7420 15108 7472
rect 15160 7460 15166 7472
rect 17218 7460 17224 7472
rect 15160 7432 17224 7460
rect 15160 7420 15166 7432
rect 17218 7420 17224 7432
rect 17276 7420 17282 7472
rect 8757 7395 8815 7401
rect 8757 7361 8769 7395
rect 8803 7361 8815 7395
rect 8757 7355 8815 7361
rect 9033 7395 9091 7401
rect 9033 7361 9045 7395
rect 9079 7392 9091 7395
rect 9674 7392 9680 7404
rect 9079 7364 9680 7392
rect 9079 7361 9091 7364
rect 9033 7355 9091 7361
rect 9674 7352 9680 7364
rect 9732 7352 9738 7404
rect 9858 7352 9864 7404
rect 9916 7352 9922 7404
rect 10137 7395 10195 7401
rect 10137 7361 10149 7395
rect 10183 7392 10195 7395
rect 10226 7392 10232 7404
rect 10183 7364 10232 7392
rect 10183 7361 10195 7364
rect 10137 7355 10195 7361
rect 10226 7352 10232 7364
rect 10284 7352 10290 7404
rect 10321 7395 10379 7401
rect 10321 7361 10333 7395
rect 10367 7361 10379 7395
rect 10321 7355 10379 7361
rect 8846 7324 8852 7336
rect 7760 7296 8852 7324
rect 8846 7284 8852 7296
rect 8904 7284 8910 7336
rect 9950 7284 9956 7336
rect 10008 7284 10014 7336
rect 2498 7216 2504 7268
rect 2556 7256 2562 7268
rect 5534 7256 5540 7268
rect 2556 7228 5540 7256
rect 2556 7216 2562 7228
rect 5534 7216 5540 7228
rect 5592 7216 5598 7268
rect 7006 7216 7012 7268
rect 7064 7256 7070 7268
rect 10336 7256 10364 7355
rect 10778 7352 10784 7404
rect 10836 7392 10842 7404
rect 10873 7395 10931 7401
rect 10873 7392 10885 7395
rect 10836 7364 10885 7392
rect 10836 7352 10842 7364
rect 10873 7361 10885 7364
rect 10919 7361 10931 7395
rect 10873 7355 10931 7361
rect 11514 7352 11520 7404
rect 11572 7352 11578 7404
rect 11606 7352 11612 7404
rect 11664 7392 11670 7404
rect 11701 7395 11759 7401
rect 11701 7392 11713 7395
rect 11664 7364 11713 7392
rect 11664 7352 11670 7364
rect 11701 7361 11713 7364
rect 11747 7361 11759 7395
rect 11701 7355 11759 7361
rect 11974 7352 11980 7404
rect 12032 7392 12038 7404
rect 14185 7395 14243 7401
rect 14185 7392 14197 7395
rect 12032 7364 14197 7392
rect 12032 7352 12038 7364
rect 14185 7361 14197 7364
rect 14231 7361 14243 7395
rect 14185 7355 14243 7361
rect 14366 7352 14372 7404
rect 14424 7352 14430 7404
rect 14458 7352 14464 7404
rect 14516 7392 14522 7404
rect 14645 7395 14703 7401
rect 14645 7392 14657 7395
rect 14516 7364 14657 7392
rect 14516 7352 14522 7364
rect 14645 7361 14657 7364
rect 14691 7361 14703 7395
rect 14645 7355 14703 7361
rect 17034 7352 17040 7404
rect 17092 7352 17098 7404
rect 10594 7284 10600 7336
rect 10652 7324 10658 7336
rect 11885 7327 11943 7333
rect 11885 7324 11897 7327
rect 10652 7296 11897 7324
rect 10652 7284 10658 7296
rect 11885 7293 11897 7296
rect 11931 7293 11943 7327
rect 12342 7324 12348 7336
rect 11885 7287 11943 7293
rect 11992 7296 12348 7324
rect 11992 7256 12020 7296
rect 12342 7284 12348 7296
rect 12400 7324 12406 7336
rect 15746 7324 15752 7336
rect 12400 7296 15752 7324
rect 12400 7284 12406 7296
rect 15746 7284 15752 7296
rect 15804 7284 15810 7336
rect 7064 7228 9076 7256
rect 10336 7228 12020 7256
rect 7064 7216 7070 7228
rect 3970 7148 3976 7200
rect 4028 7188 4034 7200
rect 8386 7188 8392 7200
rect 4028 7160 8392 7188
rect 4028 7148 4034 7160
rect 8386 7148 8392 7160
rect 8444 7148 8450 7200
rect 9048 7188 9076 7228
rect 12986 7216 12992 7268
rect 13044 7256 13050 7268
rect 13722 7256 13728 7268
rect 13044 7228 13728 7256
rect 13044 7216 13050 7228
rect 13722 7216 13728 7228
rect 13780 7216 13786 7268
rect 13906 7216 13912 7268
rect 13964 7256 13970 7268
rect 17954 7256 17960 7268
rect 13964 7228 17960 7256
rect 13964 7216 13970 7228
rect 17954 7216 17960 7228
rect 18012 7216 18018 7268
rect 10594 7188 10600 7200
rect 9048 7160 10600 7188
rect 10594 7148 10600 7160
rect 10652 7188 10658 7200
rect 11057 7191 11115 7197
rect 11057 7188 11069 7191
rect 10652 7160 11069 7188
rect 10652 7148 10658 7160
rect 11057 7157 11069 7160
rect 11103 7188 11115 7191
rect 11146 7188 11152 7200
rect 11103 7160 11152 7188
rect 11103 7157 11115 7160
rect 11057 7151 11115 7157
rect 11146 7148 11152 7160
rect 11204 7148 11210 7200
rect 11330 7148 11336 7200
rect 11388 7188 11394 7200
rect 12250 7188 12256 7200
rect 11388 7160 12256 7188
rect 11388 7148 11394 7160
rect 12250 7148 12256 7160
rect 12308 7188 12314 7200
rect 17129 7191 17187 7197
rect 17129 7188 17141 7191
rect 12308 7160 17141 7188
rect 12308 7148 12314 7160
rect 17129 7157 17141 7160
rect 17175 7157 17187 7191
rect 17129 7151 17187 7157
rect 1104 7098 18860 7120
rect 1104 7046 1950 7098
rect 2002 7046 2014 7098
rect 2066 7046 2078 7098
rect 2130 7046 2142 7098
rect 2194 7046 2206 7098
rect 2258 7046 6950 7098
rect 7002 7046 7014 7098
rect 7066 7046 7078 7098
rect 7130 7046 7142 7098
rect 7194 7046 7206 7098
rect 7258 7046 11950 7098
rect 12002 7046 12014 7098
rect 12066 7046 12078 7098
rect 12130 7046 12142 7098
rect 12194 7046 12206 7098
rect 12258 7046 16950 7098
rect 17002 7046 17014 7098
rect 17066 7046 17078 7098
rect 17130 7046 17142 7098
rect 17194 7046 17206 7098
rect 17258 7046 18860 7098
rect 1104 7024 18860 7046
rect 106 6944 112 6996
rect 164 6984 170 6996
rect 1762 6984 1768 6996
rect 164 6956 1768 6984
rect 164 6944 170 6956
rect 1762 6944 1768 6956
rect 1820 6944 1826 6996
rect 2498 6944 2504 6996
rect 2556 6984 2562 6996
rect 3142 6984 3148 6996
rect 2556 6956 3148 6984
rect 2556 6944 2562 6956
rect 3142 6944 3148 6956
rect 3200 6944 3206 6996
rect 3418 6944 3424 6996
rect 3476 6984 3482 6996
rect 4062 6984 4068 6996
rect 3476 6956 4068 6984
rect 3476 6944 3482 6956
rect 4062 6944 4068 6956
rect 4120 6944 4126 6996
rect 4338 6944 4344 6996
rect 4396 6944 4402 6996
rect 5718 6984 5724 6996
rect 4448 6956 5724 6984
rect 3878 6876 3884 6928
rect 3936 6916 3942 6928
rect 4356 6916 4384 6944
rect 3936 6888 4384 6916
rect 3936 6876 3942 6888
rect 1673 6851 1731 6857
rect 1673 6817 1685 6851
rect 1719 6848 1731 6851
rect 2314 6848 2320 6860
rect 1719 6820 2320 6848
rect 1719 6817 1731 6820
rect 1673 6811 1731 6817
rect 2314 6808 2320 6820
rect 2372 6808 2378 6860
rect 3602 6808 3608 6860
rect 3660 6808 3666 6860
rect 4338 6808 4344 6860
rect 4396 6848 4402 6860
rect 4448 6848 4476 6956
rect 5718 6944 5724 6956
rect 5776 6944 5782 6996
rect 7837 6987 7895 6993
rect 7837 6953 7849 6987
rect 7883 6984 7895 6987
rect 8018 6984 8024 6996
rect 7883 6956 8024 6984
rect 7883 6953 7895 6956
rect 7837 6947 7895 6953
rect 8018 6944 8024 6956
rect 8076 6944 8082 6996
rect 8110 6944 8116 6996
rect 8168 6984 8174 6996
rect 8754 6984 8760 6996
rect 8168 6956 8760 6984
rect 8168 6944 8174 6956
rect 8754 6944 8760 6956
rect 8812 6944 8818 6996
rect 15838 6984 15844 6996
rect 8864 6956 15844 6984
rect 5810 6916 5816 6928
rect 4540 6888 5816 6916
rect 4540 6857 4568 6888
rect 5810 6876 5816 6888
rect 5868 6876 5874 6928
rect 6454 6876 6460 6928
rect 6512 6916 6518 6928
rect 8294 6916 8300 6928
rect 6512 6888 8300 6916
rect 6512 6876 6518 6888
rect 8294 6876 8300 6888
rect 8352 6876 8358 6928
rect 8386 6876 8392 6928
rect 8444 6916 8450 6928
rect 8864 6916 8892 6956
rect 15838 6944 15844 6956
rect 15896 6944 15902 6996
rect 8444 6888 8892 6916
rect 8444 6876 8450 6888
rect 8938 6876 8944 6928
rect 8996 6916 9002 6928
rect 12897 6919 12955 6925
rect 12897 6916 12909 6919
rect 8996 6888 12909 6916
rect 8996 6876 9002 6888
rect 12897 6885 12909 6888
rect 12943 6885 12955 6919
rect 12897 6879 12955 6885
rect 4396 6820 4476 6848
rect 4525 6851 4583 6857
rect 4396 6808 4402 6820
rect 4525 6817 4537 6851
rect 4571 6817 4583 6851
rect 4525 6811 4583 6817
rect 5077 6851 5135 6857
rect 5077 6817 5089 6851
rect 5123 6848 5135 6851
rect 6086 6848 6092 6860
rect 5123 6820 6092 6848
rect 5123 6817 5135 6820
rect 5077 6811 5135 6817
rect 6086 6808 6092 6820
rect 6144 6808 6150 6860
rect 7668 6820 8340 6848
rect 1486 6672 1492 6724
rect 1544 6672 1550 6724
rect 3142 6672 3148 6724
rect 3200 6712 3206 6724
rect 3326 6712 3332 6724
rect 3200 6684 3332 6712
rect 3200 6672 3206 6684
rect 3326 6672 3332 6684
rect 3384 6672 3390 6724
rect 3620 6712 3648 6808
rect 7564 6792 7616 6798
rect 7668 6792 7696 6820
rect 3786 6740 3792 6792
rect 3844 6780 3850 6792
rect 3881 6783 3939 6789
rect 3881 6780 3893 6783
rect 3844 6752 3893 6780
rect 3844 6740 3850 6752
rect 3881 6749 3893 6752
rect 3927 6749 3939 6783
rect 3881 6743 3939 6749
rect 4062 6740 4068 6792
rect 4120 6740 4126 6792
rect 4430 6740 4436 6792
rect 4488 6740 4494 6792
rect 6638 6740 6644 6792
rect 6696 6740 6702 6792
rect 7650 6740 7656 6792
rect 7708 6740 7714 6792
rect 8018 6780 8024 6792
rect 7760 6752 8024 6780
rect 7564 6734 7616 6740
rect 3620 6684 3832 6712
rect 3804 6656 3832 6684
rect 4798 6672 4804 6724
rect 4856 6712 4862 6724
rect 5810 6712 5816 6724
rect 4856 6684 5816 6712
rect 4856 6672 4862 6684
rect 5810 6672 5816 6684
rect 5868 6712 5874 6724
rect 5868 6684 7512 6712
rect 5868 6672 5874 6684
rect 3786 6604 3792 6656
rect 3844 6604 3850 6656
rect 5074 6604 5080 6656
rect 5132 6644 5138 6656
rect 7190 6644 7196 6656
rect 5132 6616 7196 6644
rect 5132 6604 5138 6616
rect 7190 6604 7196 6616
rect 7248 6604 7254 6656
rect 7484 6644 7512 6684
rect 7760 6644 7788 6752
rect 8018 6740 8024 6752
rect 8076 6740 8082 6792
rect 8110 6740 8116 6792
rect 8168 6740 8174 6792
rect 8202 6740 8208 6792
rect 8260 6740 8266 6792
rect 8312 6656 8340 6820
rect 8846 6808 8852 6860
rect 8904 6808 8910 6860
rect 9490 6808 9496 6860
rect 9548 6848 9554 6860
rect 12802 6848 12808 6860
rect 9548 6820 12808 6848
rect 9548 6808 9554 6820
rect 12802 6808 12808 6820
rect 12860 6808 12866 6860
rect 8386 6740 8392 6792
rect 8444 6740 8450 6792
rect 8864 6780 8892 6808
rect 10870 6780 10876 6792
rect 8864 6752 10876 6780
rect 10870 6740 10876 6752
rect 10928 6740 10934 6792
rect 11054 6740 11060 6792
rect 11112 6780 11118 6792
rect 11606 6780 11612 6792
rect 11112 6752 11612 6780
rect 11112 6740 11118 6752
rect 11606 6740 11612 6752
rect 11664 6780 11670 6792
rect 12526 6780 12532 6792
rect 11664 6752 12532 6780
rect 11664 6740 11670 6752
rect 12526 6740 12532 6752
rect 12584 6740 12590 6792
rect 12618 6740 12624 6792
rect 12676 6740 12682 6792
rect 12912 6780 12940 6879
rect 13538 6876 13544 6928
rect 13596 6916 13602 6928
rect 14826 6916 14832 6928
rect 13596 6888 14832 6916
rect 13596 6876 13602 6888
rect 14826 6876 14832 6888
rect 14884 6876 14890 6928
rect 12986 6808 12992 6860
rect 13044 6848 13050 6860
rect 19242 6848 19248 6860
rect 13044 6820 19248 6848
rect 13044 6808 13050 6820
rect 19242 6808 19248 6820
rect 19300 6808 19306 6860
rect 17494 6780 17500 6792
rect 12912 6752 17500 6780
rect 17494 6740 17500 6752
rect 17552 6740 17558 6792
rect 18233 6783 18291 6789
rect 18233 6749 18245 6783
rect 18279 6780 18291 6783
rect 19426 6780 19432 6792
rect 18279 6752 19432 6780
rect 18279 6749 18291 6752
rect 18233 6743 18291 6749
rect 19426 6740 19432 6752
rect 19484 6740 19490 6792
rect 8404 6712 8432 6740
rect 12250 6712 12256 6724
rect 8404 6684 12256 6712
rect 12250 6672 12256 6684
rect 12308 6672 12314 6724
rect 16850 6712 16856 6724
rect 13004 6684 16856 6712
rect 7484 6616 7788 6644
rect 7926 6604 7932 6656
rect 7984 6644 7990 6656
rect 8202 6644 8208 6656
rect 7984 6616 8208 6644
rect 7984 6604 7990 6616
rect 8202 6604 8208 6616
rect 8260 6604 8266 6656
rect 8294 6604 8300 6656
rect 8352 6604 8358 6656
rect 8754 6604 8760 6656
rect 8812 6644 8818 6656
rect 9674 6644 9680 6656
rect 8812 6616 9680 6644
rect 8812 6604 8818 6616
rect 9674 6604 9680 6616
rect 9732 6604 9738 6656
rect 10778 6604 10784 6656
rect 10836 6644 10842 6656
rect 12526 6644 12532 6656
rect 10836 6616 12532 6644
rect 10836 6604 10842 6616
rect 12526 6604 12532 6616
rect 12584 6604 12590 6656
rect 12802 6604 12808 6656
rect 12860 6644 12866 6656
rect 13004 6644 13032 6684
rect 16850 6672 16856 6684
rect 16908 6672 16914 6724
rect 12860 6616 13032 6644
rect 13081 6647 13139 6653
rect 12860 6604 12866 6616
rect 13081 6613 13093 6647
rect 13127 6644 13139 6647
rect 13998 6644 14004 6656
rect 13127 6616 14004 6644
rect 13127 6613 13139 6616
rect 13081 6607 13139 6613
rect 13998 6604 14004 6616
rect 14056 6644 14062 6656
rect 14734 6644 14740 6656
rect 14056 6616 14740 6644
rect 14056 6604 14062 6616
rect 14734 6604 14740 6616
rect 14792 6604 14798 6656
rect 18414 6604 18420 6656
rect 18472 6604 18478 6656
rect 1104 6554 18860 6576
rect 1104 6502 2610 6554
rect 2662 6502 2674 6554
rect 2726 6502 2738 6554
rect 2790 6502 2802 6554
rect 2854 6502 2866 6554
rect 2918 6502 7610 6554
rect 7662 6502 7674 6554
rect 7726 6502 7738 6554
rect 7790 6502 7802 6554
rect 7854 6502 7866 6554
rect 7918 6502 12610 6554
rect 12662 6502 12674 6554
rect 12726 6502 12738 6554
rect 12790 6502 12802 6554
rect 12854 6502 12866 6554
rect 12918 6502 17610 6554
rect 17662 6502 17674 6554
rect 17726 6502 17738 6554
rect 17790 6502 17802 6554
rect 17854 6502 17866 6554
rect 17918 6502 18860 6554
rect 1104 6480 18860 6502
rect 4246 6449 4252 6452
rect 4233 6443 4252 6449
rect 4233 6409 4245 6443
rect 4233 6403 4252 6409
rect 4246 6400 4252 6403
rect 4304 6400 4310 6452
rect 5534 6400 5540 6452
rect 5592 6440 5598 6452
rect 7558 6440 7564 6452
rect 5592 6412 7564 6440
rect 5592 6400 5598 6412
rect 7558 6400 7564 6412
rect 7616 6400 7622 6452
rect 7926 6440 7932 6452
rect 7852 6412 7932 6440
rect 2866 6332 2872 6384
rect 2924 6372 2930 6384
rect 3142 6372 3148 6384
rect 2924 6344 3148 6372
rect 2924 6332 2930 6344
rect 3142 6332 3148 6344
rect 3200 6332 3206 6384
rect 3326 6332 3332 6384
rect 3384 6372 3390 6384
rect 3421 6375 3479 6381
rect 3421 6372 3433 6375
rect 3384 6344 3433 6372
rect 3384 6332 3390 6344
rect 3421 6341 3433 6344
rect 3467 6341 3479 6375
rect 3421 6335 3479 6341
rect 3510 6332 3516 6384
rect 3568 6372 3574 6384
rect 3568 6344 4384 6372
rect 3568 6332 3574 6344
rect 3602 6264 3608 6316
rect 3660 6264 3666 6316
rect 3712 6313 3740 6344
rect 3697 6307 3755 6313
rect 3697 6273 3709 6307
rect 3743 6273 3755 6307
rect 3697 6267 3755 6273
rect 3881 6307 3939 6313
rect 3881 6273 3893 6307
rect 3927 6273 3939 6307
rect 3881 6267 3939 6273
rect 3142 6196 3148 6248
rect 3200 6236 3206 6248
rect 3896 6236 3924 6267
rect 3970 6264 3976 6316
rect 4028 6264 4034 6316
rect 3200 6208 3924 6236
rect 3200 6196 3206 6208
rect 566 6128 572 6180
rect 624 6168 630 6180
rect 2590 6168 2596 6180
rect 624 6140 2596 6168
rect 624 6128 630 6140
rect 2590 6128 2596 6140
rect 2648 6128 2654 6180
rect 3970 6168 3976 6180
rect 2700 6140 3976 6168
rect 1578 6060 1584 6112
rect 1636 6100 1642 6112
rect 2700 6100 2728 6140
rect 3970 6128 3976 6140
rect 4028 6168 4034 6180
rect 4065 6171 4123 6177
rect 4065 6168 4077 6171
rect 4028 6140 4077 6168
rect 4028 6128 4034 6140
rect 4065 6137 4077 6140
rect 4111 6137 4123 6171
rect 4356 6168 4384 6344
rect 4430 6332 4436 6384
rect 4488 6372 4494 6384
rect 4890 6372 4896 6384
rect 4488 6344 4896 6372
rect 4488 6332 4494 6344
rect 4890 6332 4896 6344
rect 4948 6332 4954 6384
rect 7650 6372 7656 6384
rect 5000 6344 7656 6372
rect 5000 6313 5028 6344
rect 7650 6332 7656 6344
rect 7708 6332 7714 6384
rect 7852 6381 7880 6412
rect 7926 6400 7932 6412
rect 7984 6440 7990 6452
rect 8110 6440 8116 6452
rect 7984 6412 8116 6440
rect 7984 6400 7990 6412
rect 8110 6400 8116 6412
rect 8168 6400 8174 6452
rect 8205 6443 8263 6449
rect 8205 6409 8217 6443
rect 8251 6440 8263 6443
rect 8570 6440 8576 6452
rect 8251 6412 8576 6440
rect 8251 6409 8263 6412
rect 8205 6403 8263 6409
rect 8570 6400 8576 6412
rect 8628 6400 8634 6452
rect 9674 6400 9680 6452
rect 9732 6440 9738 6452
rect 9769 6443 9827 6449
rect 9769 6440 9781 6443
rect 9732 6412 9781 6440
rect 9732 6400 9738 6412
rect 9769 6409 9781 6412
rect 9815 6440 9827 6443
rect 11698 6440 11704 6452
rect 9815 6412 11704 6440
rect 9815 6409 9827 6412
rect 9769 6403 9827 6409
rect 11698 6400 11704 6412
rect 11756 6400 11762 6452
rect 12345 6443 12403 6449
rect 12345 6409 12357 6443
rect 12391 6440 12403 6443
rect 14090 6440 14096 6452
rect 12391 6412 14096 6440
rect 12391 6409 12403 6412
rect 12345 6403 12403 6409
rect 14090 6400 14096 6412
rect 14148 6400 14154 6452
rect 15930 6400 15936 6452
rect 15988 6440 15994 6452
rect 17586 6440 17592 6452
rect 15988 6412 17592 6440
rect 15988 6400 15994 6412
rect 17586 6400 17592 6412
rect 17644 6400 17650 6452
rect 7837 6375 7895 6381
rect 7837 6341 7849 6375
rect 7883 6341 7895 6375
rect 9861 6375 9919 6381
rect 9861 6372 9873 6375
rect 7837 6335 7895 6341
rect 8036 6344 9873 6372
rect 4801 6307 4859 6313
rect 4801 6273 4813 6307
rect 4847 6273 4859 6307
rect 4801 6267 4859 6273
rect 4985 6307 5043 6313
rect 4985 6273 4997 6307
rect 5031 6273 5043 6307
rect 4985 6267 5043 6273
rect 4430 6196 4436 6248
rect 4488 6236 4494 6248
rect 4816 6236 4844 6267
rect 5074 6264 5080 6316
rect 5132 6304 5138 6316
rect 5261 6307 5319 6313
rect 5261 6304 5273 6307
rect 5132 6276 5273 6304
rect 5132 6264 5138 6276
rect 5261 6273 5273 6276
rect 5307 6273 5319 6307
rect 5261 6267 5319 6273
rect 5537 6307 5595 6313
rect 5537 6273 5549 6307
rect 5583 6273 5595 6307
rect 5537 6267 5595 6273
rect 4488 6208 4844 6236
rect 5552 6236 5580 6267
rect 5718 6264 5724 6316
rect 5776 6264 5782 6316
rect 6178 6264 6184 6316
rect 6236 6304 6242 6316
rect 6638 6304 6644 6316
rect 6236 6276 6644 6304
rect 6236 6264 6242 6276
rect 6638 6264 6644 6276
rect 6696 6264 6702 6316
rect 7282 6264 7288 6316
rect 7340 6304 7346 6316
rect 8036 6313 8064 6344
rect 9861 6341 9873 6344
rect 9907 6341 9919 6375
rect 9861 6335 9919 6341
rect 10042 6332 10048 6384
rect 10100 6372 10106 6384
rect 10226 6372 10232 6384
rect 10100 6344 10232 6372
rect 10100 6332 10106 6344
rect 10226 6332 10232 6344
rect 10284 6332 10290 6384
rect 10962 6332 10968 6384
rect 11020 6372 11026 6384
rect 11790 6372 11796 6384
rect 11020 6344 11796 6372
rect 11020 6332 11026 6344
rect 11790 6332 11796 6344
rect 11848 6332 11854 6384
rect 15470 6372 15476 6384
rect 12176 6344 15476 6372
rect 8021 6307 8079 6313
rect 8021 6304 8033 6307
rect 7340 6276 8033 6304
rect 7340 6264 7346 6276
rect 8021 6273 8033 6276
rect 8067 6273 8079 6307
rect 8021 6267 8079 6273
rect 8110 6264 8116 6316
rect 8168 6264 8174 6316
rect 8202 6264 8208 6316
rect 8260 6304 8266 6316
rect 8260 6276 9628 6304
rect 8260 6264 8266 6276
rect 7098 6236 7104 6248
rect 5552 6208 7104 6236
rect 4488 6196 4494 6208
rect 7098 6196 7104 6208
rect 7156 6196 7162 6248
rect 7558 6196 7564 6248
rect 7616 6236 7622 6248
rect 8389 6239 8447 6245
rect 7616 6208 8156 6236
rect 7616 6196 7622 6208
rect 8128 6180 8156 6208
rect 8389 6205 8401 6239
rect 8435 6236 8447 6239
rect 8435 6208 8616 6236
rect 8435 6205 8447 6208
rect 8389 6199 8447 6205
rect 5534 6168 5540 6180
rect 4356 6140 5540 6168
rect 4065 6131 4123 6137
rect 5534 6128 5540 6140
rect 5592 6128 5598 6180
rect 8110 6128 8116 6180
rect 8168 6128 8174 6180
rect 8588 6168 8616 6208
rect 9490 6196 9496 6248
rect 9548 6196 9554 6248
rect 9600 6236 9628 6276
rect 9674 6264 9680 6316
rect 9732 6304 9738 6316
rect 10686 6304 10692 6316
rect 9732 6276 10692 6304
rect 9732 6264 9738 6276
rect 10686 6264 10692 6276
rect 10744 6264 10750 6316
rect 10778 6264 10784 6316
rect 10836 6304 10842 6316
rect 12176 6313 12204 6344
rect 15470 6332 15476 6344
rect 15528 6332 15534 6384
rect 12161 6307 12219 6313
rect 12161 6304 12173 6307
rect 10836 6276 12173 6304
rect 10836 6264 10842 6276
rect 12161 6273 12173 6276
rect 12207 6273 12219 6307
rect 12161 6267 12219 6273
rect 12250 6264 12256 6316
rect 12308 6304 12314 6316
rect 12345 6307 12403 6313
rect 12345 6304 12357 6307
rect 12308 6276 12357 6304
rect 12308 6264 12314 6276
rect 12345 6273 12357 6276
rect 12391 6273 12403 6307
rect 12345 6267 12403 6273
rect 13354 6264 13360 6316
rect 13412 6304 13418 6316
rect 17954 6304 17960 6316
rect 13412 6276 17960 6304
rect 13412 6264 13418 6276
rect 17954 6264 17960 6276
rect 18012 6264 18018 6316
rect 12434 6236 12440 6248
rect 9600 6208 12440 6236
rect 12434 6196 12440 6208
rect 12492 6196 12498 6248
rect 14642 6196 14648 6248
rect 14700 6196 14706 6248
rect 14660 6168 14688 6196
rect 8588 6140 14688 6168
rect 14918 6128 14924 6180
rect 14976 6168 14982 6180
rect 15746 6168 15752 6180
rect 14976 6140 15752 6168
rect 14976 6128 14982 6140
rect 15746 6128 15752 6140
rect 15804 6128 15810 6180
rect 1636 6072 2728 6100
rect 1636 6060 1642 6072
rect 3510 6060 3516 6112
rect 3568 6100 3574 6112
rect 4249 6103 4307 6109
rect 4249 6100 4261 6103
rect 3568 6072 4261 6100
rect 3568 6060 3574 6072
rect 4249 6069 4261 6072
rect 4295 6069 4307 6103
rect 4249 6063 4307 6069
rect 4614 6060 4620 6112
rect 4672 6100 4678 6112
rect 4893 6103 4951 6109
rect 4893 6100 4905 6103
rect 4672 6072 4905 6100
rect 4672 6060 4678 6072
rect 4893 6069 4905 6072
rect 4939 6100 4951 6103
rect 4982 6100 4988 6112
rect 4939 6072 4988 6100
rect 4939 6069 4951 6072
rect 4893 6063 4951 6069
rect 4982 6060 4988 6072
rect 5040 6060 5046 6112
rect 5629 6103 5687 6109
rect 5629 6069 5641 6103
rect 5675 6100 5687 6103
rect 6270 6100 6276 6112
rect 5675 6072 6276 6100
rect 5675 6069 5687 6072
rect 5629 6063 5687 6069
rect 6270 6060 6276 6072
rect 6328 6060 6334 6112
rect 7650 6060 7656 6112
rect 7708 6100 7714 6112
rect 8938 6100 8944 6112
rect 7708 6072 8944 6100
rect 7708 6060 7714 6072
rect 8938 6060 8944 6072
rect 8996 6060 9002 6112
rect 11238 6060 11244 6112
rect 11296 6100 11302 6112
rect 14458 6100 14464 6112
rect 11296 6072 14464 6100
rect 11296 6060 11302 6072
rect 14458 6060 14464 6072
rect 14516 6060 14522 6112
rect 14642 6060 14648 6112
rect 14700 6100 14706 6112
rect 16574 6100 16580 6112
rect 14700 6072 16580 6100
rect 14700 6060 14706 6072
rect 16574 6060 16580 6072
rect 16632 6060 16638 6112
rect 1104 6010 18860 6032
rect 1104 5958 1950 6010
rect 2002 5958 2014 6010
rect 2066 5958 2078 6010
rect 2130 5958 2142 6010
rect 2194 5958 2206 6010
rect 2258 5958 6950 6010
rect 7002 5958 7014 6010
rect 7066 5958 7078 6010
rect 7130 5958 7142 6010
rect 7194 5958 7206 6010
rect 7258 5958 11950 6010
rect 12002 5958 12014 6010
rect 12066 5958 12078 6010
rect 12130 5958 12142 6010
rect 12194 5958 12206 6010
rect 12258 5958 16950 6010
rect 17002 5958 17014 6010
rect 17066 5958 17078 6010
rect 17130 5958 17142 6010
rect 17194 5958 17206 6010
rect 17258 5958 18860 6010
rect 1104 5936 18860 5958
rect 2498 5856 2504 5908
rect 2556 5896 2562 5908
rect 2593 5899 2651 5905
rect 2593 5896 2605 5899
rect 2556 5868 2605 5896
rect 2556 5856 2562 5868
rect 2593 5865 2605 5868
rect 2639 5865 2651 5899
rect 2593 5859 2651 5865
rect 2682 5856 2688 5908
rect 2740 5896 2746 5908
rect 3326 5896 3332 5908
rect 2740 5868 3332 5896
rect 2740 5856 2746 5868
rect 3326 5856 3332 5868
rect 3384 5856 3390 5908
rect 3602 5856 3608 5908
rect 3660 5896 3666 5908
rect 6273 5899 6331 5905
rect 6273 5896 6285 5899
rect 3660 5868 6285 5896
rect 3660 5856 3666 5868
rect 6273 5865 6285 5868
rect 6319 5865 6331 5899
rect 6273 5859 6331 5865
rect 6380 5868 6592 5896
rect 1394 5788 1400 5840
rect 1452 5828 1458 5840
rect 6380 5828 6408 5868
rect 1452 5800 6408 5828
rect 6564 5828 6592 5868
rect 7834 5856 7840 5908
rect 7892 5896 7898 5908
rect 8846 5896 8852 5908
rect 7892 5868 8852 5896
rect 7892 5856 7898 5868
rect 8846 5856 8852 5868
rect 8904 5856 8910 5908
rect 8938 5856 8944 5908
rect 8996 5856 9002 5908
rect 10134 5896 10140 5908
rect 9048 5868 10140 5896
rect 7469 5831 7527 5837
rect 6564 5800 6868 5828
rect 1452 5788 1458 5800
rect 6840 5772 6868 5800
rect 7469 5797 7481 5831
rect 7515 5828 7527 5831
rect 9048 5828 9076 5868
rect 10134 5856 10140 5868
rect 10192 5856 10198 5908
rect 10502 5856 10508 5908
rect 10560 5856 10566 5908
rect 10870 5856 10876 5908
rect 10928 5896 10934 5908
rect 12437 5899 12495 5905
rect 12437 5896 12449 5899
rect 10928 5868 12449 5896
rect 10928 5856 10934 5868
rect 12437 5865 12449 5868
rect 12483 5865 12495 5899
rect 12437 5859 12495 5865
rect 12618 5856 12624 5908
rect 12676 5896 12682 5908
rect 12676 5868 15240 5896
rect 12676 5856 12682 5868
rect 7515 5800 9076 5828
rect 7515 5797 7527 5800
rect 7469 5791 7527 5797
rect 9122 5788 9128 5840
rect 9180 5828 9186 5840
rect 11057 5831 11115 5837
rect 11057 5828 11069 5831
rect 9180 5800 11069 5828
rect 9180 5788 9186 5800
rect 11057 5797 11069 5800
rect 11103 5797 11115 5831
rect 15102 5828 15108 5840
rect 11057 5791 11115 5797
rect 11532 5800 13814 5828
rect 842 5720 848 5772
rect 900 5760 906 5772
rect 2685 5763 2743 5769
rect 2685 5760 2697 5763
rect 900 5732 2697 5760
rect 900 5720 906 5732
rect 2685 5729 2697 5732
rect 2731 5760 2743 5763
rect 2866 5760 2872 5772
rect 2731 5732 2872 5760
rect 2731 5729 2743 5732
rect 2685 5723 2743 5729
rect 2866 5720 2872 5732
rect 2924 5720 2930 5772
rect 3053 5763 3111 5769
rect 3053 5729 3065 5763
rect 3099 5760 3111 5763
rect 3418 5760 3424 5772
rect 3099 5732 3424 5760
rect 3099 5729 3111 5732
rect 3053 5723 3111 5729
rect 2406 5652 2412 5704
rect 2464 5652 2470 5704
rect 2501 5695 2559 5701
rect 2501 5661 2513 5695
rect 2547 5692 2559 5695
rect 2590 5692 2596 5704
rect 2547 5664 2596 5692
rect 2547 5661 2559 5664
rect 2501 5655 2559 5661
rect 2590 5652 2596 5664
rect 2648 5652 2654 5704
rect 750 5584 756 5636
rect 808 5624 814 5636
rect 808 5596 2268 5624
rect 808 5584 814 5596
rect 1302 5516 1308 5568
rect 1360 5556 1366 5568
rect 1486 5556 1492 5568
rect 1360 5528 1492 5556
rect 1360 5516 1366 5528
rect 1486 5516 1492 5528
rect 1544 5516 1550 5568
rect 2240 5556 2268 5596
rect 2314 5584 2320 5636
rect 2372 5624 2378 5636
rect 3068 5624 3096 5723
rect 3418 5720 3424 5732
rect 3476 5720 3482 5772
rect 3881 5763 3939 5769
rect 3881 5729 3893 5763
rect 3927 5760 3939 5763
rect 4062 5760 4068 5772
rect 3927 5732 4068 5760
rect 3927 5729 3939 5732
rect 3881 5723 3939 5729
rect 4062 5720 4068 5732
rect 4120 5720 4126 5772
rect 4341 5763 4399 5769
rect 4341 5729 4353 5763
rect 4387 5760 4399 5763
rect 4798 5760 4804 5772
rect 4387 5732 4804 5760
rect 4387 5729 4399 5732
rect 4341 5723 4399 5729
rect 4798 5720 4804 5732
rect 4856 5720 4862 5772
rect 4890 5720 4896 5772
rect 4948 5760 4954 5772
rect 5994 5760 6000 5772
rect 4948 5732 6000 5760
rect 4948 5720 4954 5732
rect 5994 5720 6000 5732
rect 6052 5720 6058 5772
rect 6638 5720 6644 5772
rect 6696 5720 6702 5772
rect 6822 5720 6828 5772
rect 6880 5720 6886 5772
rect 11532 5760 11560 5800
rect 9048 5732 11560 5760
rect 11609 5763 11667 5769
rect 4157 5695 4215 5701
rect 4157 5661 4169 5695
rect 4203 5692 4215 5695
rect 4522 5692 4528 5704
rect 4203 5664 4528 5692
rect 4203 5661 4215 5664
rect 4157 5655 4215 5661
rect 4522 5652 4528 5664
rect 4580 5652 4586 5704
rect 6454 5652 6460 5704
rect 6512 5692 6518 5704
rect 6549 5695 6607 5701
rect 6549 5692 6561 5695
rect 6512 5664 6561 5692
rect 6512 5652 6518 5664
rect 6549 5661 6561 5664
rect 6595 5661 6607 5695
rect 6549 5655 6607 5661
rect 7466 5652 7472 5704
rect 7524 5652 7530 5704
rect 7650 5652 7656 5704
rect 7708 5692 7714 5704
rect 7745 5695 7803 5701
rect 7745 5692 7757 5695
rect 7708 5664 7757 5692
rect 7708 5652 7714 5664
rect 7745 5661 7757 5664
rect 7791 5661 7803 5695
rect 7745 5655 7803 5661
rect 8294 5652 8300 5704
rect 8352 5692 8358 5704
rect 8938 5692 8944 5704
rect 8352 5664 8944 5692
rect 8352 5652 8358 5664
rect 8938 5652 8944 5664
rect 8996 5692 9002 5704
rect 9048 5692 9076 5732
rect 8996 5664 9076 5692
rect 8996 5652 9002 5664
rect 9122 5652 9128 5704
rect 9180 5652 9186 5704
rect 3789 5627 3847 5633
rect 3789 5624 3801 5627
rect 2372 5596 3096 5624
rect 3252 5596 3801 5624
rect 2372 5584 2378 5596
rect 3252 5556 3280 5596
rect 3789 5593 3801 5596
rect 3835 5593 3847 5627
rect 3789 5587 3847 5593
rect 4172 5596 8340 5624
rect 4172 5568 4200 5596
rect 2240 5528 3280 5556
rect 3513 5559 3571 5565
rect 3513 5525 3525 5559
rect 3559 5556 3571 5559
rect 3602 5556 3608 5568
rect 3559 5528 3608 5556
rect 3559 5525 3571 5528
rect 3513 5519 3571 5525
rect 3602 5516 3608 5528
rect 3660 5516 3666 5568
rect 4154 5516 4160 5568
rect 4212 5516 4218 5568
rect 5258 5516 5264 5568
rect 5316 5556 5322 5568
rect 5810 5556 5816 5568
rect 5316 5528 5816 5556
rect 5316 5516 5322 5528
rect 5810 5516 5816 5528
rect 5868 5516 5874 5568
rect 6730 5516 6736 5568
rect 6788 5556 6794 5568
rect 7834 5556 7840 5568
rect 6788 5528 7840 5556
rect 6788 5516 6794 5528
rect 7834 5516 7840 5528
rect 7892 5516 7898 5568
rect 7926 5516 7932 5568
rect 7984 5556 7990 5568
rect 8202 5556 8208 5568
rect 7984 5528 8208 5556
rect 7984 5516 7990 5528
rect 8202 5516 8208 5528
rect 8260 5516 8266 5568
rect 8312 5556 8340 5596
rect 8386 5584 8392 5636
rect 8444 5624 8450 5636
rect 9324 5633 9352 5732
rect 11609 5729 11621 5763
rect 11655 5760 11667 5763
rect 13538 5760 13544 5772
rect 11655 5732 13544 5760
rect 11655 5729 11667 5732
rect 11609 5723 11667 5729
rect 13538 5720 13544 5732
rect 13596 5720 13602 5772
rect 9493 5695 9551 5701
rect 9493 5661 9505 5695
rect 9539 5692 9551 5695
rect 9950 5692 9956 5704
rect 9539 5664 9956 5692
rect 9539 5661 9551 5664
rect 9493 5655 9551 5661
rect 9950 5652 9956 5664
rect 10008 5652 10014 5704
rect 10505 5695 10563 5701
rect 10505 5661 10517 5695
rect 10551 5692 10563 5695
rect 10594 5692 10600 5704
rect 10551 5664 10600 5692
rect 10551 5661 10563 5664
rect 10505 5655 10563 5661
rect 10594 5652 10600 5664
rect 10652 5652 10658 5704
rect 10781 5695 10839 5701
rect 10781 5661 10793 5695
rect 10827 5661 10839 5695
rect 10781 5655 10839 5661
rect 9217 5627 9275 5633
rect 9217 5624 9229 5627
rect 8444 5596 9229 5624
rect 8444 5584 8450 5596
rect 9217 5593 9229 5596
rect 9263 5593 9275 5627
rect 9217 5587 9275 5593
rect 9309 5627 9367 5633
rect 9309 5593 9321 5627
rect 9355 5593 9367 5627
rect 9309 5587 9367 5593
rect 9766 5584 9772 5636
rect 9824 5624 9830 5636
rect 10689 5627 10747 5633
rect 10689 5624 10701 5627
rect 9824 5596 10701 5624
rect 9824 5584 9830 5596
rect 10612 5568 10640 5596
rect 10689 5593 10701 5596
rect 10735 5593 10747 5627
rect 10796 5624 10824 5655
rect 11146 5652 11152 5704
rect 11204 5692 11210 5704
rect 11241 5695 11299 5701
rect 11241 5692 11253 5695
rect 11204 5664 11253 5692
rect 11204 5652 11210 5664
rect 11241 5661 11253 5664
rect 11287 5661 11299 5695
rect 11241 5655 11299 5661
rect 11333 5695 11391 5701
rect 11333 5661 11345 5695
rect 11379 5692 11391 5695
rect 11698 5692 11704 5704
rect 11379 5664 11704 5692
rect 11379 5661 11391 5664
rect 11333 5655 11391 5661
rect 11698 5652 11704 5664
rect 11756 5652 11762 5704
rect 11790 5652 11796 5704
rect 11848 5652 11854 5704
rect 12529 5695 12587 5701
rect 12529 5661 12541 5695
rect 12575 5692 12587 5695
rect 13170 5692 13176 5704
rect 12575 5664 13176 5692
rect 12575 5661 12587 5664
rect 12529 5655 12587 5661
rect 13170 5652 13176 5664
rect 13228 5652 13234 5704
rect 13786 5692 13814 5800
rect 14384 5800 15108 5828
rect 13998 5720 14004 5772
rect 14056 5760 14062 5772
rect 14384 5769 14412 5800
rect 15102 5788 15108 5800
rect 15160 5788 15166 5840
rect 15212 5828 15240 5868
rect 16850 5856 16856 5908
rect 16908 5896 16914 5908
rect 17221 5899 17279 5905
rect 17221 5896 17233 5899
rect 16908 5868 17233 5896
rect 16908 5856 16914 5868
rect 17221 5865 17233 5868
rect 17267 5865 17279 5899
rect 17221 5859 17279 5865
rect 16022 5828 16028 5840
rect 15212 5800 16028 5828
rect 16022 5788 16028 5800
rect 16080 5788 16086 5840
rect 14369 5763 14427 5769
rect 14369 5760 14381 5763
rect 14056 5732 14381 5760
rect 14056 5720 14062 5732
rect 14369 5729 14381 5732
rect 14415 5729 14427 5763
rect 14369 5723 14427 5729
rect 14458 5720 14464 5772
rect 14516 5720 14522 5772
rect 14826 5720 14832 5772
rect 14884 5760 14890 5772
rect 16482 5760 16488 5772
rect 14884 5732 16488 5760
rect 14884 5720 14890 5732
rect 16482 5720 16488 5732
rect 16540 5720 16546 5772
rect 16574 5720 16580 5772
rect 16632 5720 16638 5772
rect 14553 5695 14611 5701
rect 14553 5692 14565 5695
rect 13786 5664 14565 5692
rect 14553 5661 14565 5664
rect 14599 5661 14611 5695
rect 14553 5655 14611 5661
rect 14645 5695 14703 5701
rect 14645 5661 14657 5695
rect 14691 5692 14703 5695
rect 15102 5692 15108 5704
rect 14691 5664 15108 5692
rect 14691 5661 14703 5664
rect 14645 5655 14703 5661
rect 14568 5624 14596 5655
rect 15102 5652 15108 5664
rect 15160 5652 15166 5704
rect 15194 5652 15200 5704
rect 15252 5652 15258 5704
rect 15565 5695 15623 5701
rect 15565 5661 15577 5695
rect 15611 5661 15623 5695
rect 15565 5655 15623 5661
rect 14918 5624 14924 5636
rect 10796 5596 12388 5624
rect 10689 5587 10747 5593
rect 9122 5556 9128 5568
rect 8312 5528 9128 5556
rect 9122 5516 9128 5528
rect 9180 5516 9186 5568
rect 10594 5516 10600 5568
rect 10652 5516 10658 5568
rect 10778 5516 10784 5568
rect 10836 5556 10842 5568
rect 11425 5559 11483 5565
rect 11425 5556 11437 5559
rect 10836 5528 11437 5556
rect 10836 5516 10842 5528
rect 11425 5525 11437 5528
rect 11471 5556 11483 5559
rect 11606 5556 11612 5568
rect 11471 5528 11612 5556
rect 11471 5525 11483 5528
rect 11425 5519 11483 5525
rect 11606 5516 11612 5528
rect 11664 5516 11670 5568
rect 12360 5556 12388 5596
rect 14117 5596 14504 5624
rect 14568 5596 14924 5624
rect 14117 5556 14145 5596
rect 12360 5528 14145 5556
rect 14182 5516 14188 5568
rect 14240 5516 14246 5568
rect 14476 5556 14504 5596
rect 14918 5584 14924 5596
rect 14976 5584 14982 5636
rect 15580 5624 15608 5655
rect 16298 5652 16304 5704
rect 16356 5692 16362 5704
rect 16669 5695 16727 5701
rect 16669 5692 16681 5695
rect 16356 5664 16681 5692
rect 16356 5652 16362 5664
rect 16669 5661 16681 5664
rect 16715 5661 16727 5695
rect 16669 5655 16727 5661
rect 16758 5652 16764 5704
rect 16816 5652 16822 5704
rect 16853 5695 16911 5701
rect 16853 5661 16865 5695
rect 16899 5661 16911 5695
rect 16853 5655 16911 5661
rect 16574 5624 16580 5636
rect 15580 5596 16580 5624
rect 16574 5584 16580 5596
rect 16632 5584 16638 5636
rect 14826 5556 14832 5568
rect 14476 5528 14832 5556
rect 14826 5516 14832 5528
rect 14884 5516 14890 5568
rect 15194 5516 15200 5568
rect 15252 5556 15258 5568
rect 16393 5559 16451 5565
rect 16393 5556 16405 5559
rect 15252 5528 16405 5556
rect 15252 5516 15258 5528
rect 16393 5525 16405 5528
rect 16439 5525 16451 5559
rect 16868 5556 16896 5655
rect 17236 5624 17264 5859
rect 17954 5856 17960 5908
rect 18012 5896 18018 5908
rect 18049 5899 18107 5905
rect 18049 5896 18061 5899
rect 18012 5868 18061 5896
rect 18012 5856 18018 5868
rect 18049 5865 18061 5868
rect 18095 5865 18107 5899
rect 18049 5859 18107 5865
rect 17310 5720 17316 5772
rect 17368 5760 17374 5772
rect 17368 5732 17908 5760
rect 17368 5720 17374 5732
rect 17586 5652 17592 5704
rect 17644 5652 17650 5704
rect 17880 5701 17908 5732
rect 17865 5695 17923 5701
rect 17865 5661 17877 5695
rect 17911 5661 17923 5695
rect 17865 5655 17923 5661
rect 17681 5627 17739 5633
rect 17681 5624 17693 5627
rect 17236 5596 17693 5624
rect 17681 5593 17693 5596
rect 17727 5593 17739 5627
rect 18322 5624 18328 5636
rect 17681 5587 17739 5593
rect 17972 5596 18328 5624
rect 17972 5556 18000 5596
rect 18322 5584 18328 5596
rect 18380 5584 18386 5636
rect 16868 5528 18000 5556
rect 16393 5519 16451 5525
rect 1104 5466 18860 5488
rect 1104 5414 2610 5466
rect 2662 5414 2674 5466
rect 2726 5414 2738 5466
rect 2790 5414 2802 5466
rect 2854 5414 2866 5466
rect 2918 5414 7610 5466
rect 7662 5414 7674 5466
rect 7726 5414 7738 5466
rect 7790 5414 7802 5466
rect 7854 5414 7866 5466
rect 7918 5414 12610 5466
rect 12662 5414 12674 5466
rect 12726 5414 12738 5466
rect 12790 5414 12802 5466
rect 12854 5414 12866 5466
rect 12918 5414 17610 5466
rect 17662 5414 17674 5466
rect 17726 5414 17738 5466
rect 17790 5414 17802 5466
rect 17854 5414 17866 5466
rect 17918 5414 18860 5466
rect 1104 5392 18860 5414
rect 1118 5312 1124 5364
rect 1176 5352 1182 5364
rect 1302 5352 1308 5364
rect 1176 5324 1308 5352
rect 1176 5312 1182 5324
rect 1302 5312 1308 5324
rect 1360 5312 1366 5364
rect 3050 5312 3056 5364
rect 3108 5352 3114 5364
rect 3108 5324 6224 5352
rect 3108 5312 3114 5324
rect 2406 5244 2412 5296
rect 2464 5284 2470 5296
rect 3418 5284 3424 5296
rect 2464 5256 3424 5284
rect 2464 5244 2470 5256
rect 3418 5244 3424 5256
rect 3476 5244 3482 5296
rect 3602 5244 3608 5296
rect 3660 5284 3666 5296
rect 5902 5284 5908 5296
rect 3660 5256 4752 5284
rect 3660 5244 3666 5256
rect 3050 5176 3056 5228
rect 3108 5216 3114 5228
rect 3145 5219 3203 5225
rect 3145 5216 3157 5219
rect 3108 5188 3157 5216
rect 3108 5176 3114 5188
rect 3145 5185 3157 5188
rect 3191 5185 3203 5219
rect 3145 5179 3203 5185
rect 3789 5219 3847 5225
rect 3789 5185 3801 5219
rect 3835 5216 3847 5219
rect 3970 5216 3976 5228
rect 3835 5188 3976 5216
rect 3835 5185 3847 5188
rect 3789 5179 3847 5185
rect 3970 5176 3976 5188
rect 4028 5176 4034 5228
rect 4154 5176 4160 5228
rect 4212 5176 4218 5228
rect 4338 5176 4344 5228
rect 4396 5216 4402 5228
rect 4724 5225 4752 5256
rect 4816 5256 5908 5284
rect 4433 5219 4491 5225
rect 4433 5216 4445 5219
rect 4396 5188 4445 5216
rect 4396 5176 4402 5188
rect 4433 5185 4445 5188
rect 4479 5185 4491 5219
rect 4433 5179 4491 5185
rect 4698 5219 4756 5225
rect 4698 5185 4710 5219
rect 4744 5185 4756 5219
rect 4698 5179 4756 5185
rect 4062 5108 4068 5160
rect 4120 5108 4126 5160
rect 4816 5148 4844 5256
rect 5902 5244 5908 5256
rect 5960 5244 5966 5296
rect 4982 5176 4988 5228
rect 5040 5176 5046 5228
rect 5166 5176 5172 5228
rect 5224 5176 5230 5228
rect 5626 5176 5632 5228
rect 5684 5176 5690 5228
rect 6196 5216 6224 5324
rect 7282 5312 7288 5364
rect 7340 5312 7346 5364
rect 7466 5312 7472 5364
rect 7524 5352 7530 5364
rect 7742 5352 7748 5364
rect 7524 5324 7748 5352
rect 7524 5312 7530 5324
rect 7742 5312 7748 5324
rect 7800 5352 7806 5364
rect 10594 5352 10600 5364
rect 7800 5324 10600 5352
rect 7800 5312 7806 5324
rect 10594 5312 10600 5324
rect 10652 5312 10658 5364
rect 10870 5312 10876 5364
rect 10928 5352 10934 5364
rect 11514 5352 11520 5364
rect 10928 5324 11520 5352
rect 10928 5312 10934 5324
rect 11514 5312 11520 5324
rect 11572 5312 11578 5364
rect 11624 5324 12664 5352
rect 6564 5256 8432 5284
rect 6365 5219 6423 5225
rect 6365 5216 6377 5219
rect 6196 5188 6377 5216
rect 6365 5185 6377 5188
rect 6411 5216 6423 5219
rect 6454 5216 6460 5228
rect 6411 5188 6460 5216
rect 6411 5185 6423 5188
rect 6365 5179 6423 5185
rect 6454 5176 6460 5188
rect 6512 5176 6518 5228
rect 6564 5225 6592 5256
rect 6549 5219 6607 5225
rect 6549 5185 6561 5219
rect 6595 5185 6607 5219
rect 6549 5179 6607 5185
rect 6917 5219 6975 5225
rect 6917 5185 6929 5219
rect 6963 5185 6975 5219
rect 6917 5179 6975 5185
rect 6564 5148 6592 5179
rect 4172 5120 4844 5148
rect 4908 5120 6592 5148
rect 4172 5092 4200 5120
rect 4154 5040 4160 5092
rect 4212 5040 4218 5092
rect 4798 5040 4804 5092
rect 4856 5040 4862 5092
rect 4338 4972 4344 5024
rect 4396 5012 4402 5024
rect 4908 5012 4936 5120
rect 5258 5040 5264 5092
rect 5316 5080 5322 5092
rect 6932 5080 6960 5179
rect 7282 5176 7288 5228
rect 7340 5216 7346 5228
rect 7653 5219 7711 5225
rect 7653 5216 7665 5219
rect 7340 5188 7665 5216
rect 7340 5176 7346 5188
rect 7653 5185 7665 5188
rect 7699 5185 7711 5219
rect 7653 5179 7711 5185
rect 7926 5176 7932 5228
rect 7984 5176 7990 5228
rect 8110 5176 8116 5228
rect 8168 5216 8174 5228
rect 8297 5219 8355 5225
rect 8297 5216 8309 5219
rect 8168 5188 8309 5216
rect 8168 5176 8174 5188
rect 8297 5185 8309 5188
rect 8343 5185 8355 5219
rect 8404 5216 8432 5256
rect 8846 5244 8852 5296
rect 8904 5244 8910 5296
rect 10410 5284 10416 5296
rect 8956 5256 10416 5284
rect 8956 5216 8984 5256
rect 10410 5244 10416 5256
rect 10468 5244 10474 5296
rect 10502 5244 10508 5296
rect 10560 5284 10566 5296
rect 11624 5284 11652 5324
rect 12526 5284 12532 5296
rect 10560 5256 11652 5284
rect 11900 5256 12532 5284
rect 10560 5244 10566 5256
rect 8404 5188 8984 5216
rect 8297 5179 8355 5185
rect 9030 5176 9036 5228
rect 9088 5176 9094 5228
rect 9122 5176 9128 5228
rect 9180 5216 9186 5228
rect 10962 5216 10968 5228
rect 9180 5188 10968 5216
rect 9180 5176 9186 5188
rect 10962 5176 10968 5188
rect 11020 5176 11026 5228
rect 11900 5225 11928 5256
rect 12526 5244 12532 5256
rect 12584 5244 12590 5296
rect 12636 5293 12664 5324
rect 16390 5312 16396 5364
rect 16448 5352 16454 5364
rect 16448 5324 16896 5352
rect 16448 5312 16454 5324
rect 12621 5287 12679 5293
rect 12621 5253 12633 5287
rect 12667 5253 12679 5287
rect 12621 5247 12679 5253
rect 16482 5244 16488 5296
rect 16540 5284 16546 5296
rect 16868 5293 16896 5324
rect 17494 5312 17500 5364
rect 17552 5312 17558 5364
rect 16669 5287 16727 5293
rect 16669 5284 16681 5287
rect 16540 5256 16681 5284
rect 16540 5244 16546 5256
rect 16669 5253 16681 5256
rect 16715 5253 16727 5287
rect 16669 5247 16727 5253
rect 16853 5287 16911 5293
rect 16853 5253 16865 5287
rect 16899 5284 16911 5287
rect 16899 5256 18552 5284
rect 16899 5253 16911 5256
rect 16853 5247 16911 5253
rect 11885 5219 11943 5225
rect 11885 5185 11897 5219
rect 11931 5185 11943 5219
rect 11885 5179 11943 5185
rect 12250 5176 12256 5228
rect 12308 5216 12314 5228
rect 12345 5219 12403 5225
rect 12345 5216 12357 5219
rect 12308 5188 12357 5216
rect 12308 5176 12314 5188
rect 12345 5185 12357 5188
rect 12391 5185 12403 5219
rect 12345 5179 12403 5185
rect 12437 5219 12495 5225
rect 12437 5185 12449 5219
rect 12483 5216 12495 5219
rect 13446 5216 13452 5228
rect 12483 5188 13452 5216
rect 12483 5185 12495 5188
rect 12437 5179 12495 5185
rect 13446 5176 13452 5188
rect 13504 5176 13510 5228
rect 15470 5176 15476 5228
rect 15528 5176 15534 5228
rect 15654 5176 15660 5228
rect 15712 5176 15718 5228
rect 17405 5219 17463 5225
rect 17405 5185 17417 5219
rect 17451 5185 17463 5219
rect 17405 5179 17463 5185
rect 17589 5219 17647 5225
rect 17589 5185 17601 5219
rect 17635 5216 17647 5219
rect 17954 5216 17960 5228
rect 17635 5188 17960 5216
rect 17635 5185 17647 5188
rect 17589 5179 17647 5185
rect 7006 5108 7012 5160
rect 7064 5108 7070 5160
rect 7466 5108 7472 5160
rect 7524 5148 7530 5160
rect 7837 5151 7895 5157
rect 7837 5148 7849 5151
rect 7524 5120 7849 5148
rect 7524 5108 7530 5120
rect 7837 5117 7849 5120
rect 7883 5117 7895 5151
rect 8938 5148 8944 5160
rect 7837 5111 7895 5117
rect 8680 5120 8944 5148
rect 8680 5092 8708 5120
rect 8938 5108 8944 5120
rect 8996 5148 9002 5160
rect 9217 5151 9275 5157
rect 9217 5148 9229 5151
rect 8996 5120 9229 5148
rect 8996 5108 9002 5120
rect 9217 5117 9229 5120
rect 9263 5117 9275 5151
rect 11701 5151 11759 5157
rect 11701 5148 11713 5151
rect 9217 5111 9275 5117
rect 9416 5120 11713 5148
rect 8386 5080 8392 5092
rect 5316 5052 6960 5080
rect 8220 5052 8392 5080
rect 5316 5040 5322 5052
rect 4396 4984 4936 5012
rect 4396 4972 4402 4984
rect 5718 4972 5724 5024
rect 5776 4972 5782 5024
rect 5994 4972 6000 5024
rect 6052 5012 6058 5024
rect 6089 5015 6147 5021
rect 6089 5012 6101 5015
rect 6052 4984 6101 5012
rect 6052 4972 6058 4984
rect 6089 4981 6101 4984
rect 6135 4981 6147 5015
rect 6089 4975 6147 4981
rect 6730 4972 6736 5024
rect 6788 5012 6794 5024
rect 8220 5012 8248 5052
rect 8386 5040 8392 5052
rect 8444 5040 8450 5092
rect 8662 5040 8668 5092
rect 8720 5040 8726 5092
rect 6788 4984 8248 5012
rect 6788 4972 6794 4984
rect 8294 4972 8300 5024
rect 8352 5012 8358 5024
rect 9416 5012 9444 5120
rect 11701 5117 11713 5120
rect 11747 5148 11759 5151
rect 11790 5148 11796 5160
rect 11747 5120 11796 5148
rect 11747 5117 11759 5120
rect 11701 5111 11759 5117
rect 11790 5108 11796 5120
rect 11848 5108 11854 5160
rect 12069 5151 12127 5157
rect 12069 5117 12081 5151
rect 12115 5148 12127 5151
rect 13078 5148 13084 5160
rect 12115 5120 13084 5148
rect 12115 5117 12127 5120
rect 12069 5111 12127 5117
rect 13078 5108 13084 5120
rect 13136 5148 13142 5160
rect 16114 5148 16120 5160
rect 13136 5120 16120 5148
rect 13136 5108 13142 5120
rect 16114 5108 16120 5120
rect 16172 5108 16178 5160
rect 16482 5108 16488 5160
rect 16540 5108 16546 5160
rect 16666 5108 16672 5160
rect 16724 5108 16730 5160
rect 16758 5108 16764 5160
rect 16816 5148 16822 5160
rect 17420 5148 17448 5179
rect 17954 5176 17960 5188
rect 18012 5176 18018 5228
rect 18322 5176 18328 5228
rect 18380 5176 18386 5228
rect 18524 5225 18552 5256
rect 18509 5219 18567 5225
rect 18509 5185 18521 5219
rect 18555 5185 18567 5219
rect 18509 5179 18567 5185
rect 16816 5120 17448 5148
rect 16816 5108 16822 5120
rect 10042 5040 10048 5092
rect 10100 5080 10106 5092
rect 16684 5080 16712 5108
rect 10100 5052 16712 5080
rect 10100 5040 10106 5052
rect 8352 4984 9444 5012
rect 8352 4972 8358 4984
rect 10594 4972 10600 5024
rect 10652 5012 10658 5024
rect 12250 5012 12256 5024
rect 10652 4984 12256 5012
rect 10652 4972 10658 4984
rect 12250 4972 12256 4984
rect 12308 4972 12314 5024
rect 12526 4972 12532 5024
rect 12584 5012 12590 5024
rect 12621 5015 12679 5021
rect 12621 5012 12633 5015
rect 12584 4984 12633 5012
rect 12584 4972 12590 4984
rect 12621 4981 12633 4984
rect 12667 4981 12679 5015
rect 12621 4975 12679 4981
rect 16666 4972 16672 5024
rect 16724 5012 16730 5024
rect 17037 5015 17095 5021
rect 17037 5012 17049 5015
rect 16724 4984 17049 5012
rect 16724 4972 16730 4984
rect 17037 4981 17049 4984
rect 17083 4981 17095 5015
rect 17037 4975 17095 4981
rect 18322 4972 18328 5024
rect 18380 4972 18386 5024
rect 1104 4922 18860 4944
rect 1104 4870 1950 4922
rect 2002 4870 2014 4922
rect 2066 4870 2078 4922
rect 2130 4870 2142 4922
rect 2194 4870 2206 4922
rect 2258 4870 6950 4922
rect 7002 4870 7014 4922
rect 7066 4870 7078 4922
rect 7130 4870 7142 4922
rect 7194 4870 7206 4922
rect 7258 4870 11950 4922
rect 12002 4870 12014 4922
rect 12066 4870 12078 4922
rect 12130 4870 12142 4922
rect 12194 4870 12206 4922
rect 12258 4870 16950 4922
rect 17002 4870 17014 4922
rect 17066 4870 17078 4922
rect 17130 4870 17142 4922
rect 17194 4870 17206 4922
rect 17258 4870 18860 4922
rect 1104 4848 18860 4870
rect 1762 4768 1768 4820
rect 1820 4808 1826 4820
rect 1946 4808 1952 4820
rect 1820 4780 1952 4808
rect 1820 4768 1826 4780
rect 1946 4768 1952 4780
rect 2004 4768 2010 4820
rect 2498 4768 2504 4820
rect 2556 4808 2562 4820
rect 5074 4808 5080 4820
rect 2556 4780 5080 4808
rect 2556 4768 2562 4780
rect 5074 4768 5080 4780
rect 5132 4768 5138 4820
rect 5261 4811 5319 4817
rect 5261 4777 5273 4811
rect 5307 4808 5319 4811
rect 5442 4808 5448 4820
rect 5307 4780 5448 4808
rect 5307 4777 5319 4780
rect 5261 4771 5319 4777
rect 5442 4768 5448 4780
rect 5500 4768 5506 4820
rect 5721 4811 5779 4817
rect 5721 4777 5733 4811
rect 5767 4808 5779 4811
rect 5810 4808 5816 4820
rect 5767 4780 5816 4808
rect 5767 4777 5779 4780
rect 5721 4771 5779 4777
rect 5810 4768 5816 4780
rect 5868 4808 5874 4820
rect 6730 4808 6736 4820
rect 5868 4780 6736 4808
rect 5868 4768 5874 4780
rect 6730 4768 6736 4780
rect 6788 4768 6794 4820
rect 7374 4808 7380 4820
rect 7111 4780 7380 4808
rect 2774 4700 2780 4752
rect 2832 4700 2838 4752
rect 4246 4740 4252 4752
rect 3160 4712 4252 4740
rect 1762 4632 1768 4684
rect 1820 4672 1826 4684
rect 1820 4644 2912 4672
rect 1820 4632 1826 4644
rect 1673 4607 1731 4613
rect 1673 4573 1685 4607
rect 1719 4573 1731 4607
rect 1673 4567 1731 4573
rect 2041 4607 2099 4613
rect 2041 4573 2053 4607
rect 2087 4573 2099 4607
rect 2041 4567 2099 4573
rect 2317 4607 2375 4613
rect 2317 4573 2329 4607
rect 2363 4604 2375 4607
rect 2406 4604 2412 4616
rect 2363 4576 2412 4604
rect 2363 4573 2375 4576
rect 2317 4567 2375 4573
rect 1688 4468 1716 4567
rect 2056 4536 2084 4567
rect 2406 4564 2412 4576
rect 2464 4564 2470 4616
rect 2884 4613 2912 4644
rect 2869 4607 2927 4613
rect 2869 4573 2881 4607
rect 2915 4604 2927 4607
rect 3160 4604 3188 4712
rect 4246 4700 4252 4712
rect 4304 4700 4310 4752
rect 5166 4700 5172 4752
rect 5224 4740 5230 4752
rect 5353 4743 5411 4749
rect 5353 4740 5365 4743
rect 5224 4712 5365 4740
rect 5224 4700 5230 4712
rect 5353 4709 5365 4712
rect 5399 4709 5411 4743
rect 7006 4740 7012 4752
rect 5353 4703 5411 4709
rect 6886 4712 7012 4740
rect 3234 4632 3240 4684
rect 3292 4672 3298 4684
rect 3881 4675 3939 4681
rect 3881 4672 3893 4675
rect 3292 4644 3893 4672
rect 3292 4632 3298 4644
rect 3881 4641 3893 4644
rect 3927 4641 3939 4675
rect 3881 4635 3939 4641
rect 4341 4675 4399 4681
rect 4341 4641 4353 4675
rect 4387 4672 4399 4675
rect 4430 4672 4436 4684
rect 4387 4644 4436 4672
rect 4387 4641 4399 4644
rect 4341 4635 4399 4641
rect 4430 4632 4436 4644
rect 4488 4632 4494 4684
rect 4706 4632 4712 4684
rect 4764 4672 4770 4684
rect 4893 4675 4951 4681
rect 4893 4672 4905 4675
rect 4764 4644 4905 4672
rect 4764 4632 4770 4644
rect 4893 4641 4905 4644
rect 4939 4641 4951 4675
rect 4893 4635 4951 4641
rect 5077 4675 5135 4681
rect 5077 4641 5089 4675
rect 5123 4672 5135 4675
rect 6886 4672 6914 4712
rect 7006 4700 7012 4712
rect 7064 4700 7070 4752
rect 7111 4681 7139 4780
rect 7374 4768 7380 4780
rect 7432 4768 7438 4820
rect 7837 4811 7895 4817
rect 7837 4777 7849 4811
rect 7883 4808 7895 4811
rect 9950 4808 9956 4820
rect 7883 4780 9956 4808
rect 7883 4777 7895 4780
rect 7837 4771 7895 4777
rect 9950 4768 9956 4780
rect 10008 4768 10014 4820
rect 11977 4811 12035 4817
rect 11977 4777 11989 4811
rect 12023 4808 12035 4811
rect 12066 4808 12072 4820
rect 12023 4780 12072 4808
rect 12023 4777 12035 4780
rect 11977 4771 12035 4777
rect 12066 4768 12072 4780
rect 12124 4768 12130 4820
rect 12176 4780 14596 4808
rect 7190 4700 7196 4752
rect 7248 4700 7254 4752
rect 7561 4743 7619 4749
rect 7561 4709 7573 4743
rect 7607 4740 7619 4743
rect 9122 4740 9128 4752
rect 7607 4712 9128 4740
rect 7607 4709 7619 4712
rect 7561 4703 7619 4709
rect 9122 4700 9128 4712
rect 9180 4700 9186 4752
rect 9674 4700 9680 4752
rect 9732 4740 9738 4752
rect 12176 4740 12204 4780
rect 14461 4743 14519 4749
rect 14461 4740 14473 4743
rect 9732 4712 12204 4740
rect 12268 4712 14473 4740
rect 9732 4700 9738 4712
rect 5123 4644 6914 4672
rect 7101 4675 7159 4681
rect 5123 4641 5135 4644
rect 5077 4635 5135 4641
rect 7101 4641 7113 4675
rect 7147 4641 7159 4675
rect 7208 4672 7236 4700
rect 12268 4672 12296 4712
rect 14461 4709 14473 4712
rect 14507 4709 14519 4743
rect 14568 4740 14596 4780
rect 14642 4768 14648 4820
rect 14700 4768 14706 4820
rect 15286 4808 15292 4820
rect 14752 4780 15292 4808
rect 14752 4740 14780 4780
rect 15286 4768 15292 4780
rect 15344 4768 15350 4820
rect 14568 4712 14780 4740
rect 14461 4703 14519 4709
rect 14826 4700 14832 4752
rect 14884 4700 14890 4752
rect 14844 4672 14872 4700
rect 15565 4675 15623 4681
rect 7208 4644 12296 4672
rect 12406 4644 14412 4672
rect 14844 4644 15240 4672
rect 7101 4635 7159 4641
rect 2915 4576 3188 4604
rect 2915 4573 2927 4576
rect 2869 4567 2927 4573
rect 3970 4564 3976 4616
rect 4028 4564 4034 4616
rect 4154 4564 4160 4616
rect 4212 4604 4218 4616
rect 4801 4607 4859 4613
rect 4801 4604 4813 4607
rect 4212 4576 4813 4604
rect 4212 4564 4218 4576
rect 4801 4573 4813 4576
rect 4847 4573 4859 4607
rect 4801 4567 4859 4573
rect 4985 4607 5043 4613
rect 4985 4573 4997 4607
rect 5031 4573 5043 4607
rect 4985 4567 5043 4573
rect 4338 4536 4344 4548
rect 2056 4508 4344 4536
rect 4338 4496 4344 4508
rect 4396 4496 4402 4548
rect 4706 4496 4712 4548
rect 4764 4536 4770 4548
rect 5000 4536 5028 4567
rect 5534 4564 5540 4616
rect 5592 4564 5598 4616
rect 5813 4607 5871 4613
rect 5813 4573 5825 4607
rect 5859 4604 5871 4607
rect 5859 4576 6776 4604
rect 5859 4573 5871 4576
rect 5813 4567 5871 4573
rect 4764 4508 5028 4536
rect 4764 4496 4770 4508
rect 6086 4468 6092 4480
rect 1688 4440 6092 4468
rect 6086 4428 6092 4440
rect 6144 4428 6150 4480
rect 6748 4468 6776 4576
rect 7190 4564 7196 4616
rect 7248 4564 7254 4616
rect 7285 4607 7343 4613
rect 7285 4573 7297 4607
rect 7331 4573 7343 4607
rect 7285 4567 7343 4573
rect 7377 4607 7435 4613
rect 7377 4573 7389 4607
rect 7423 4573 7435 4607
rect 7377 4567 7435 4573
rect 7641 4607 7699 4613
rect 7641 4573 7653 4607
rect 7687 4604 7699 4607
rect 7742 4604 7748 4616
rect 7687 4576 7748 4604
rect 7687 4573 7699 4576
rect 7641 4567 7699 4573
rect 6822 4496 6828 4548
rect 6880 4536 6886 4548
rect 7300 4536 7328 4567
rect 6880 4508 7328 4536
rect 7392 4536 7420 4567
rect 7742 4564 7748 4576
rect 7800 4564 7806 4616
rect 7837 4607 7895 4613
rect 7837 4573 7849 4607
rect 7883 4604 7895 4607
rect 8018 4604 8024 4616
rect 7883 4576 8024 4604
rect 7883 4573 7895 4576
rect 7837 4567 7895 4573
rect 8018 4564 8024 4576
rect 8076 4564 8082 4616
rect 8110 4564 8116 4616
rect 8168 4604 8174 4616
rect 8570 4604 8576 4616
rect 8168 4576 8576 4604
rect 8168 4564 8174 4576
rect 8570 4564 8576 4576
rect 8628 4564 8634 4616
rect 10410 4564 10416 4616
rect 10468 4564 10474 4616
rect 10686 4564 10692 4616
rect 10744 4604 10750 4616
rect 11241 4607 11299 4613
rect 11241 4604 11253 4607
rect 10744 4576 11253 4604
rect 10744 4564 10750 4576
rect 11241 4573 11253 4576
rect 11287 4573 11299 4607
rect 11241 4567 11299 4573
rect 11514 4564 11520 4616
rect 11572 4564 11578 4616
rect 11790 4564 11796 4616
rect 11848 4564 11854 4616
rect 11882 4564 11888 4616
rect 11940 4604 11946 4616
rect 12406 4604 12434 4644
rect 11940 4576 12434 4604
rect 11940 4564 11946 4576
rect 13538 4564 13544 4616
rect 13596 4604 13602 4616
rect 14277 4607 14335 4613
rect 14277 4604 14289 4607
rect 13596 4576 14289 4604
rect 13596 4564 13602 4576
rect 14277 4573 14289 4576
rect 14323 4573 14335 4607
rect 14277 4567 14335 4573
rect 8846 4536 8852 4548
rect 7392 4508 8852 4536
rect 6880 4496 6886 4508
rect 8846 4496 8852 4508
rect 8904 4496 8910 4548
rect 9950 4496 9956 4548
rect 10008 4536 10014 4548
rect 13262 4536 13268 4548
rect 10008 4508 13268 4536
rect 10008 4496 10014 4508
rect 13262 4496 13268 4508
rect 13320 4496 13326 4548
rect 14384 4545 14412 4644
rect 14550 4564 14556 4616
rect 14608 4564 14614 4616
rect 14642 4564 14648 4616
rect 14700 4564 14706 4616
rect 14734 4564 14740 4616
rect 14792 4604 14798 4616
rect 14829 4607 14887 4613
rect 14829 4604 14841 4607
rect 14792 4576 14841 4604
rect 14792 4564 14798 4576
rect 14829 4573 14841 4576
rect 14875 4573 14887 4607
rect 14829 4567 14887 4573
rect 15010 4564 15016 4616
rect 15068 4564 15074 4616
rect 15212 4613 15240 4644
rect 15565 4641 15577 4675
rect 15611 4672 15623 4675
rect 15930 4672 15936 4684
rect 15611 4644 15936 4672
rect 15611 4641 15623 4644
rect 15565 4635 15623 4641
rect 15930 4632 15936 4644
rect 15988 4632 15994 4684
rect 15197 4607 15255 4613
rect 15197 4573 15209 4607
rect 15243 4604 15255 4607
rect 16114 4604 16120 4616
rect 15243 4576 16120 4604
rect 15243 4573 15255 4576
rect 15197 4567 15255 4573
rect 16114 4564 16120 4576
rect 16172 4604 16178 4616
rect 16298 4604 16304 4616
rect 16172 4576 16304 4604
rect 16172 4564 16178 4576
rect 16298 4564 16304 4576
rect 16356 4564 16362 4616
rect 14369 4539 14427 4545
rect 14369 4505 14381 4539
rect 14415 4505 14427 4539
rect 14369 4499 14427 4505
rect 8754 4468 8760 4480
rect 6748 4440 8760 4468
rect 8754 4428 8760 4440
rect 8812 4428 8818 4480
rect 10686 4428 10692 4480
rect 10744 4468 10750 4480
rect 11609 4471 11667 4477
rect 11609 4468 11621 4471
rect 10744 4440 11621 4468
rect 10744 4428 10750 4440
rect 11609 4437 11621 4440
rect 11655 4468 11667 4471
rect 18966 4468 18972 4480
rect 11655 4440 18972 4468
rect 11655 4437 11667 4440
rect 11609 4431 11667 4437
rect 18966 4428 18972 4440
rect 19024 4428 19030 4480
rect 1104 4378 18860 4400
rect 1104 4326 2610 4378
rect 2662 4326 2674 4378
rect 2726 4326 2738 4378
rect 2790 4326 2802 4378
rect 2854 4326 2866 4378
rect 2918 4326 7610 4378
rect 7662 4326 7674 4378
rect 7726 4326 7738 4378
rect 7790 4326 7802 4378
rect 7854 4326 7866 4378
rect 7918 4326 12610 4378
rect 12662 4326 12674 4378
rect 12726 4326 12738 4378
rect 12790 4326 12802 4378
rect 12854 4326 12866 4378
rect 12918 4326 17610 4378
rect 17662 4326 17674 4378
rect 17726 4326 17738 4378
rect 17790 4326 17802 4378
rect 17854 4326 17866 4378
rect 17918 4326 18860 4378
rect 1104 4304 18860 4326
rect 2317 4267 2375 4273
rect 2317 4233 2329 4267
rect 2363 4264 2375 4267
rect 2363 4236 2452 4264
rect 2363 4233 2375 4236
rect 2317 4227 2375 4233
rect 1854 4156 1860 4208
rect 1912 4196 1918 4208
rect 2424 4196 2452 4236
rect 2590 4224 2596 4276
rect 2648 4264 2654 4276
rect 3878 4264 3884 4276
rect 2648 4236 3884 4264
rect 2648 4224 2654 4236
rect 3878 4224 3884 4236
rect 3936 4224 3942 4276
rect 4430 4224 4436 4276
rect 4488 4264 4494 4276
rect 5074 4264 5080 4276
rect 4488 4236 5080 4264
rect 4488 4224 4494 4236
rect 5074 4224 5080 4236
rect 5132 4224 5138 4276
rect 5166 4224 5172 4276
rect 5224 4264 5230 4276
rect 5629 4267 5687 4273
rect 5224 4236 5488 4264
rect 5224 4224 5230 4236
rect 5460 4196 5488 4236
rect 5629 4233 5641 4267
rect 5675 4264 5687 4267
rect 12986 4264 12992 4276
rect 5675 4236 12992 4264
rect 5675 4233 5687 4236
rect 5629 4227 5687 4233
rect 12986 4224 12992 4236
rect 13044 4264 13050 4276
rect 15194 4264 15200 4276
rect 13044 4236 15200 4264
rect 13044 4224 13050 4236
rect 15194 4224 15200 4236
rect 15252 4224 15258 4276
rect 5810 4196 5816 4208
rect 1912 4168 2360 4196
rect 2424 4168 3280 4196
rect 1912 4156 1918 4168
rect 1670 4088 1676 4140
rect 1728 4128 1734 4140
rect 2041 4131 2099 4137
rect 1728 4100 1992 4128
rect 1728 4088 1734 4100
rect 1857 4063 1915 4069
rect 1857 4029 1869 4063
rect 1903 4029 1915 4063
rect 1964 4060 1992 4100
rect 2041 4097 2053 4131
rect 2087 4128 2099 4131
rect 2222 4128 2228 4140
rect 2087 4100 2228 4128
rect 2087 4097 2099 4100
rect 2041 4091 2099 4097
rect 2222 4088 2228 4100
rect 2280 4088 2286 4140
rect 2332 4128 2360 4168
rect 2685 4131 2743 4137
rect 2685 4128 2697 4131
rect 2332 4100 2697 4128
rect 2685 4097 2697 4100
rect 2731 4097 2743 4131
rect 2685 4091 2743 4097
rect 2409 4063 2467 4069
rect 2409 4060 2421 4063
rect 1964 4032 2421 4060
rect 1857 4023 1915 4029
rect 2409 4029 2421 4032
rect 2455 4029 2467 4063
rect 2409 4023 2467 4029
rect 2501 4063 2559 4069
rect 2501 4029 2513 4063
rect 2547 4029 2559 4063
rect 3252 4060 3280 4168
rect 3344 4168 5396 4196
rect 5460 4168 5816 4196
rect 3344 4137 3372 4168
rect 3329 4131 3387 4137
rect 3329 4097 3341 4131
rect 3375 4097 3387 4131
rect 3329 4091 3387 4097
rect 3697 4131 3755 4137
rect 3697 4097 3709 4131
rect 3743 4128 3755 4131
rect 3878 4128 3884 4140
rect 3743 4100 3884 4128
rect 3743 4097 3755 4100
rect 3697 4091 3755 4097
rect 3878 4088 3884 4100
rect 3936 4088 3942 4140
rect 3973 4131 4031 4137
rect 3973 4097 3985 4131
rect 4019 4128 4031 4131
rect 4246 4128 4252 4140
rect 4019 4100 4252 4128
rect 4019 4097 4031 4100
rect 3973 4091 4031 4097
rect 4246 4088 4252 4100
rect 4304 4088 4310 4140
rect 4338 4088 4344 4140
rect 4396 4088 4402 4140
rect 4614 4088 4620 4140
rect 4672 4088 4678 4140
rect 5258 4088 5264 4140
rect 5316 4088 5322 4140
rect 5368 4128 5396 4168
rect 5810 4156 5816 4168
rect 5868 4156 5874 4208
rect 6454 4156 6460 4208
rect 6512 4196 6518 4208
rect 6512 4168 8156 4196
rect 6512 4156 6518 4168
rect 7466 4128 7472 4140
rect 5368 4100 7472 4128
rect 7466 4088 7472 4100
rect 7524 4088 7530 4140
rect 8128 4128 8156 4168
rect 8294 4156 8300 4208
rect 8352 4196 8358 4208
rect 8481 4199 8539 4205
rect 8481 4196 8493 4199
rect 8352 4168 8493 4196
rect 8352 4156 8358 4168
rect 8481 4165 8493 4168
rect 8527 4165 8539 4199
rect 8481 4159 8539 4165
rect 8754 4156 8760 4208
rect 8812 4196 8818 4208
rect 9398 4196 9404 4208
rect 8812 4168 9404 4196
rect 8812 4156 8818 4168
rect 9398 4156 9404 4168
rect 9456 4156 9462 4208
rect 9950 4156 9956 4208
rect 10008 4196 10014 4208
rect 11974 4196 11980 4208
rect 10008 4168 11980 4196
rect 10008 4156 10014 4168
rect 11974 4156 11980 4168
rect 12032 4196 12038 4208
rect 13078 4196 13084 4208
rect 12032 4168 12204 4196
rect 12032 4156 12038 4168
rect 9125 4131 9183 4137
rect 9125 4128 9137 4131
rect 8128 4100 9137 4128
rect 9125 4097 9137 4100
rect 9171 4097 9183 4131
rect 9677 4131 9735 4137
rect 9677 4128 9689 4131
rect 9125 4091 9183 4097
rect 9232 4100 9689 4128
rect 4798 4060 4804 4072
rect 3252 4032 4804 4060
rect 2501 4023 2559 4029
rect 1872 3924 1900 4023
rect 2314 3952 2320 4004
rect 2372 3992 2378 4004
rect 2516 3992 2544 4023
rect 4798 4020 4804 4032
rect 4856 4020 4862 4072
rect 5169 4063 5227 4069
rect 5169 4029 5181 4063
rect 5215 4060 5227 4063
rect 5442 4060 5448 4072
rect 5215 4032 5448 4060
rect 5215 4029 5227 4032
rect 5169 4023 5227 4029
rect 5442 4020 5448 4032
rect 5500 4020 5506 4072
rect 5534 4020 5540 4072
rect 5592 4060 5598 4072
rect 9232 4060 9260 4100
rect 9677 4097 9689 4100
rect 9723 4097 9735 4131
rect 9677 4091 9735 4097
rect 9861 4131 9919 4137
rect 9861 4097 9873 4131
rect 9907 4128 9919 4131
rect 10962 4128 10968 4140
rect 9907 4100 10968 4128
rect 9907 4097 9919 4100
rect 9861 4091 9919 4097
rect 10962 4088 10968 4100
rect 11020 4088 11026 4140
rect 11146 4088 11152 4140
rect 11204 4128 11210 4140
rect 12176 4137 12204 4168
rect 12452 4168 13084 4196
rect 12069 4131 12127 4137
rect 12069 4128 12081 4131
rect 11204 4100 12081 4128
rect 11204 4088 11210 4100
rect 12069 4097 12081 4100
rect 12115 4097 12127 4131
rect 12069 4091 12127 4097
rect 12161 4131 12219 4137
rect 12161 4097 12173 4131
rect 12207 4097 12219 4131
rect 12161 4091 12219 4097
rect 12253 4131 12311 4137
rect 12253 4097 12265 4131
rect 12299 4128 12311 4131
rect 12342 4128 12348 4140
rect 12299 4100 12348 4128
rect 12299 4097 12311 4100
rect 12253 4091 12311 4097
rect 12342 4088 12348 4100
rect 12400 4088 12406 4140
rect 12452 4137 12480 4168
rect 13078 4156 13084 4168
rect 13136 4156 13142 4208
rect 16390 4156 16396 4208
rect 16448 4196 16454 4208
rect 16761 4199 16819 4205
rect 16761 4196 16773 4199
rect 16448 4168 16773 4196
rect 16448 4156 16454 4168
rect 16761 4165 16773 4168
rect 16807 4165 16819 4199
rect 16761 4159 16819 4165
rect 12437 4131 12495 4137
rect 12437 4097 12449 4131
rect 12483 4097 12495 4131
rect 12437 4091 12495 4097
rect 12621 4131 12679 4137
rect 12621 4097 12633 4131
rect 12667 4128 12679 4131
rect 13906 4128 13912 4140
rect 12667 4100 13912 4128
rect 12667 4097 12679 4100
rect 12621 4091 12679 4097
rect 13906 4088 13912 4100
rect 13964 4088 13970 4140
rect 14918 4088 14924 4140
rect 14976 4128 14982 4140
rect 17310 4128 17316 4140
rect 14976 4100 17316 4128
rect 14976 4088 14982 4100
rect 17310 4088 17316 4100
rect 17368 4088 17374 4140
rect 18230 4088 18236 4140
rect 18288 4088 18294 4140
rect 5592 4032 9260 4060
rect 5592 4020 5598 4032
rect 9582 4020 9588 4072
rect 9640 4020 9646 4072
rect 9766 4020 9772 4072
rect 9824 4020 9830 4072
rect 10042 4020 10048 4072
rect 10100 4020 10106 4072
rect 10410 4020 10416 4072
rect 10468 4060 10474 4072
rect 11330 4060 11336 4072
rect 10468 4032 11336 4060
rect 10468 4020 10474 4032
rect 11330 4020 11336 4032
rect 11388 4020 11394 4072
rect 11790 4020 11796 4072
rect 11848 4060 11854 4072
rect 11977 4063 12035 4069
rect 11977 4060 11989 4063
rect 11848 4032 11989 4060
rect 11848 4020 11854 4032
rect 11977 4029 11989 4032
rect 12023 4029 12035 4063
rect 11977 4023 12035 4029
rect 12529 4063 12587 4069
rect 12529 4029 12541 4063
rect 12575 4060 12587 4063
rect 12575 4032 13584 4060
rect 12575 4029 12587 4032
rect 12529 4023 12587 4029
rect 2372 3964 2544 3992
rect 2372 3952 2378 3964
rect 4338 3952 4344 4004
rect 4396 3992 4402 4004
rect 13446 3992 13452 4004
rect 4396 3964 13452 3992
rect 4396 3952 4402 3964
rect 13446 3952 13452 3964
rect 13504 3952 13510 4004
rect 13556 3992 13584 4032
rect 13722 4020 13728 4072
rect 13780 4060 13786 4072
rect 17954 4060 17960 4072
rect 13780 4032 17960 4060
rect 13780 4020 13786 4032
rect 17954 4020 17960 4032
rect 18012 4020 18018 4072
rect 13556 3964 14228 3992
rect 2958 3924 2964 3936
rect 1872 3896 2964 3924
rect 2958 3884 2964 3896
rect 3016 3924 3022 3936
rect 4890 3924 4896 3936
rect 3016 3896 4896 3924
rect 3016 3884 3022 3896
rect 4890 3884 4896 3896
rect 4948 3884 4954 3936
rect 5442 3884 5448 3936
rect 5500 3884 5506 3936
rect 5629 3927 5687 3933
rect 5629 3893 5641 3927
rect 5675 3924 5687 3927
rect 5902 3924 5908 3936
rect 5675 3896 5908 3924
rect 5675 3893 5687 3896
rect 5629 3887 5687 3893
rect 5902 3884 5908 3896
rect 5960 3884 5966 3936
rect 6454 3884 6460 3936
rect 6512 3924 6518 3936
rect 8294 3924 8300 3936
rect 6512 3896 8300 3924
rect 6512 3884 6518 3896
rect 8294 3884 8300 3896
rect 8352 3884 8358 3936
rect 9398 3884 9404 3936
rect 9456 3924 9462 3936
rect 11146 3924 11152 3936
rect 9456 3896 11152 3924
rect 9456 3884 9462 3896
rect 11146 3884 11152 3896
rect 11204 3884 11210 3936
rect 11514 3884 11520 3936
rect 11572 3924 11578 3936
rect 11793 3927 11851 3933
rect 11793 3924 11805 3927
rect 11572 3896 11805 3924
rect 11572 3884 11578 3896
rect 11793 3893 11805 3896
rect 11839 3893 11851 3927
rect 14200 3924 14228 3964
rect 14366 3952 14372 4004
rect 14424 3992 14430 4004
rect 14918 3992 14924 4004
rect 14424 3964 14924 3992
rect 14424 3952 14430 3964
rect 14918 3952 14924 3964
rect 14976 3952 14982 4004
rect 15102 3952 15108 4004
rect 15160 3992 15166 4004
rect 17862 3992 17868 4004
rect 15160 3964 17868 3992
rect 15160 3952 15166 3964
rect 17862 3952 17868 3964
rect 17920 3952 17926 4004
rect 15378 3924 15384 3936
rect 14200 3896 15384 3924
rect 11793 3887 11851 3893
rect 15378 3884 15384 3896
rect 15436 3884 15442 3936
rect 16853 3927 16911 3933
rect 16853 3893 16865 3927
rect 16899 3924 16911 3927
rect 17402 3924 17408 3936
rect 16899 3896 17408 3924
rect 16899 3893 16911 3896
rect 16853 3887 16911 3893
rect 17402 3884 17408 3896
rect 17460 3884 17466 3936
rect 18414 3884 18420 3936
rect 18472 3884 18478 3936
rect 1104 3834 18860 3856
rect 1104 3782 1950 3834
rect 2002 3782 2014 3834
rect 2066 3782 2078 3834
rect 2130 3782 2142 3834
rect 2194 3782 2206 3834
rect 2258 3782 6950 3834
rect 7002 3782 7014 3834
rect 7066 3782 7078 3834
rect 7130 3782 7142 3834
rect 7194 3782 7206 3834
rect 7258 3782 11950 3834
rect 12002 3782 12014 3834
rect 12066 3782 12078 3834
rect 12130 3782 12142 3834
rect 12194 3782 12206 3834
rect 12258 3782 16950 3834
rect 17002 3782 17014 3834
rect 17066 3782 17078 3834
rect 17130 3782 17142 3834
rect 17194 3782 17206 3834
rect 17258 3782 18860 3834
rect 1104 3760 18860 3782
rect 290 3680 296 3732
rect 348 3720 354 3732
rect 5442 3720 5448 3732
rect 348 3692 5448 3720
rect 348 3680 354 3692
rect 5442 3680 5448 3692
rect 5500 3680 5506 3732
rect 6362 3720 6368 3732
rect 5552 3692 6368 3720
rect 1026 3612 1032 3664
rect 1084 3652 1090 3664
rect 2314 3652 2320 3664
rect 1084 3624 2320 3652
rect 1084 3612 1090 3624
rect 2314 3612 2320 3624
rect 2372 3612 2378 3664
rect 3050 3612 3056 3664
rect 3108 3652 3114 3664
rect 5552 3652 5580 3692
rect 6362 3680 6368 3692
rect 6420 3680 6426 3732
rect 6917 3723 6975 3729
rect 6917 3689 6929 3723
rect 6963 3720 6975 3723
rect 9674 3720 9680 3732
rect 6963 3692 9680 3720
rect 6963 3689 6975 3692
rect 6917 3683 6975 3689
rect 9674 3680 9680 3692
rect 9732 3680 9738 3732
rect 10226 3680 10232 3732
rect 10284 3720 10290 3732
rect 11422 3720 11428 3732
rect 10284 3692 11428 3720
rect 10284 3680 10290 3692
rect 11422 3680 11428 3692
rect 11480 3680 11486 3732
rect 11698 3680 11704 3732
rect 11756 3720 11762 3732
rect 16390 3720 16396 3732
rect 11756 3692 16396 3720
rect 11756 3680 11762 3692
rect 16390 3680 16396 3692
rect 16448 3680 16454 3732
rect 16574 3680 16580 3732
rect 16632 3720 16638 3732
rect 17129 3723 17187 3729
rect 17129 3720 17141 3723
rect 16632 3692 17141 3720
rect 16632 3680 16638 3692
rect 17129 3689 17141 3692
rect 17175 3689 17187 3723
rect 17129 3683 17187 3689
rect 17862 3680 17868 3732
rect 17920 3680 17926 3732
rect 17954 3680 17960 3732
rect 18012 3720 18018 3732
rect 18049 3723 18107 3729
rect 18049 3720 18061 3723
rect 18012 3692 18061 3720
rect 18012 3680 18018 3692
rect 18049 3689 18061 3692
rect 18095 3689 18107 3723
rect 18049 3683 18107 3689
rect 3108 3624 5580 3652
rect 3108 3612 3114 3624
rect 5626 3612 5632 3664
rect 5684 3652 5690 3664
rect 8941 3655 8999 3661
rect 8941 3652 8953 3655
rect 5684 3624 8953 3652
rect 5684 3612 5690 3624
rect 8941 3621 8953 3624
rect 8987 3621 8999 3655
rect 10870 3652 10876 3664
rect 8941 3615 8999 3621
rect 9600 3624 10876 3652
rect 1673 3587 1731 3593
rect 1673 3553 1685 3587
rect 1719 3584 1731 3587
rect 2866 3584 2872 3596
rect 1719 3556 2872 3584
rect 1719 3553 1731 3556
rect 1673 3547 1731 3553
rect 2866 3544 2872 3556
rect 2924 3544 2930 3596
rect 5810 3544 5816 3596
rect 5868 3584 5874 3596
rect 6546 3584 6552 3596
rect 5868 3556 6552 3584
rect 5868 3544 5874 3556
rect 6546 3544 6552 3556
rect 6604 3544 6610 3596
rect 7282 3584 7288 3596
rect 7208 3556 7288 3584
rect 4617 3529 4675 3535
rect 1394 3476 1400 3528
rect 1452 3476 1458 3528
rect 1854 3476 1860 3528
rect 1912 3516 1918 3528
rect 2041 3519 2099 3525
rect 2041 3516 2053 3519
rect 1912 3488 2053 3516
rect 1912 3476 1918 3488
rect 2041 3485 2053 3488
rect 2087 3485 2099 3519
rect 2041 3479 2099 3485
rect 2682 3476 2688 3528
rect 2740 3476 2746 3528
rect 2777 3519 2835 3525
rect 2777 3485 2789 3519
rect 2823 3485 2835 3519
rect 2777 3479 2835 3485
rect 1394 3340 1400 3392
rect 1452 3380 1458 3392
rect 1946 3380 1952 3392
rect 1452 3352 1952 3380
rect 1452 3340 1458 3352
rect 1946 3340 1952 3352
rect 2004 3340 2010 3392
rect 2501 3383 2559 3389
rect 2501 3349 2513 3383
rect 2547 3380 2559 3383
rect 2792 3380 2820 3479
rect 3050 3476 3056 3528
rect 3108 3476 3114 3528
rect 4154 3476 4160 3528
rect 4212 3476 4218 3528
rect 4338 3476 4344 3528
rect 4396 3476 4402 3528
rect 4522 3476 4528 3528
rect 4580 3476 4586 3528
rect 4617 3495 4629 3529
rect 4663 3516 4675 3529
rect 5258 3516 5264 3528
rect 4663 3495 5264 3516
rect 4617 3489 5264 3495
rect 4632 3488 5264 3489
rect 5258 3476 5264 3488
rect 5316 3476 5322 3528
rect 5997 3519 6055 3525
rect 5997 3516 6009 3519
rect 5368 3488 6009 3516
rect 3234 3408 3240 3460
rect 3292 3448 3298 3460
rect 4249 3451 4307 3457
rect 3292 3420 4108 3448
rect 3292 3408 3298 3420
rect 2547 3352 2820 3380
rect 2547 3349 2559 3352
rect 2501 3343 2559 3349
rect 2958 3340 2964 3392
rect 3016 3380 3022 3392
rect 3973 3383 4031 3389
rect 3973 3380 3985 3383
rect 3016 3352 3985 3380
rect 3016 3340 3022 3352
rect 3973 3349 3985 3352
rect 4019 3349 4031 3383
rect 4080 3380 4108 3420
rect 4249 3417 4261 3451
rect 4295 3448 4307 3451
rect 4890 3448 4896 3460
rect 4295 3420 4896 3448
rect 4295 3417 4307 3420
rect 4249 3411 4307 3417
rect 4890 3408 4896 3420
rect 4948 3408 4954 3460
rect 5368 3380 5396 3488
rect 5997 3485 6009 3488
rect 6043 3516 6055 3519
rect 6086 3516 6092 3528
rect 6043 3488 6092 3516
rect 6043 3485 6055 3488
rect 5997 3479 6055 3485
rect 6086 3476 6092 3488
rect 6144 3476 6150 3528
rect 6181 3519 6239 3525
rect 6181 3485 6193 3519
rect 6227 3516 6239 3519
rect 6914 3516 6920 3528
rect 6227 3488 6920 3516
rect 6227 3485 6239 3488
rect 6181 3479 6239 3485
rect 5534 3408 5540 3460
rect 5592 3448 5598 3460
rect 6196 3448 6224 3479
rect 6914 3476 6920 3488
rect 6972 3476 6978 3528
rect 7006 3476 7012 3528
rect 7064 3525 7070 3528
rect 7208 3525 7236 3556
rect 7282 3544 7288 3556
rect 7340 3544 7346 3596
rect 8110 3584 8116 3596
rect 7484 3556 8116 3584
rect 7064 3519 7107 3525
rect 7095 3485 7107 3519
rect 7064 3479 7107 3485
rect 7193 3519 7251 3525
rect 7193 3485 7205 3519
rect 7239 3485 7251 3519
rect 7193 3479 7251 3485
rect 7064 3476 7070 3479
rect 7374 3476 7380 3528
rect 7432 3516 7438 3528
rect 7484 3525 7512 3556
rect 8110 3544 8116 3556
rect 8168 3544 8174 3596
rect 9600 3584 9628 3624
rect 10870 3612 10876 3624
rect 10928 3612 10934 3664
rect 12802 3652 12808 3664
rect 11716 3624 12808 3652
rect 8588 3556 9628 3584
rect 7469 3519 7527 3525
rect 7469 3516 7481 3519
rect 7432 3488 7481 3516
rect 7432 3476 7438 3488
rect 7469 3485 7481 3488
rect 7515 3485 7527 3519
rect 7469 3479 7527 3485
rect 7929 3519 7987 3525
rect 7929 3485 7941 3519
rect 7975 3485 7987 3519
rect 7929 3479 7987 3485
rect 5592 3420 6224 3448
rect 5592 3408 5598 3420
rect 6362 3408 6368 3460
rect 6420 3408 6426 3460
rect 7285 3451 7343 3457
rect 7285 3417 7297 3451
rect 7331 3448 7343 3451
rect 7944 3448 7972 3479
rect 8202 3476 8208 3528
rect 8260 3476 8266 3528
rect 8294 3476 8300 3528
rect 8352 3476 8358 3528
rect 8588 3525 8616 3556
rect 9674 3544 9680 3596
rect 9732 3584 9738 3596
rect 11716 3584 11744 3624
rect 12802 3612 12808 3624
rect 12860 3612 12866 3664
rect 12897 3655 12955 3661
rect 12897 3621 12909 3655
rect 12943 3652 12955 3655
rect 13170 3652 13176 3664
rect 12943 3624 13176 3652
rect 12943 3621 12955 3624
rect 12897 3615 12955 3621
rect 13170 3612 13176 3624
rect 13228 3652 13234 3664
rect 13228 3624 17264 3652
rect 13228 3612 13234 3624
rect 9732 3556 11744 3584
rect 9732 3544 9738 3556
rect 11790 3544 11796 3596
rect 11848 3584 11854 3596
rect 13998 3584 14004 3596
rect 11848 3556 14004 3584
rect 11848 3544 11854 3556
rect 13998 3544 14004 3556
rect 14056 3544 14062 3596
rect 15286 3544 15292 3596
rect 15344 3584 15350 3596
rect 15746 3584 15752 3596
rect 15344 3556 15752 3584
rect 15344 3544 15350 3556
rect 15746 3544 15752 3556
rect 15804 3544 15810 3596
rect 15930 3544 15936 3596
rect 15988 3544 15994 3596
rect 16132 3556 17080 3584
rect 8573 3519 8631 3525
rect 8573 3485 8585 3519
rect 8619 3485 8631 3519
rect 9125 3519 9183 3525
rect 8573 3479 8631 3485
rect 8680 3488 9076 3516
rect 8478 3448 8484 3460
rect 7331 3420 7880 3448
rect 7944 3420 8484 3448
rect 7331 3417 7343 3420
rect 7285 3411 7343 3417
rect 4080 3352 5396 3380
rect 3973 3343 4031 3349
rect 5626 3340 5632 3392
rect 5684 3380 5690 3392
rect 7745 3383 7803 3389
rect 7745 3380 7757 3383
rect 5684 3352 7757 3380
rect 5684 3340 5690 3352
rect 7745 3349 7757 3352
rect 7791 3349 7803 3383
rect 7852 3380 7880 3420
rect 8478 3408 8484 3420
rect 8536 3448 8542 3460
rect 8680 3448 8708 3488
rect 8536 3420 8708 3448
rect 8536 3408 8542 3420
rect 8754 3408 8760 3460
rect 8812 3408 8818 3460
rect 9048 3448 9076 3488
rect 9125 3485 9137 3519
rect 9171 3516 9183 3519
rect 9214 3516 9220 3528
rect 9171 3488 9220 3516
rect 9171 3485 9183 3488
rect 9125 3479 9183 3485
rect 9214 3476 9220 3488
rect 9272 3476 9278 3528
rect 9306 3476 9312 3528
rect 9364 3476 9370 3528
rect 9401 3519 9459 3525
rect 9401 3485 9413 3519
rect 9447 3516 9459 3519
rect 9490 3516 9496 3528
rect 9447 3488 9496 3516
rect 9447 3485 9459 3488
rect 9401 3479 9459 3485
rect 9490 3476 9496 3488
rect 9548 3476 9554 3528
rect 11882 3516 11888 3528
rect 9600 3488 11888 3516
rect 9600 3448 9628 3488
rect 11882 3476 11888 3488
rect 11940 3476 11946 3528
rect 12618 3476 12624 3528
rect 12676 3476 12682 3528
rect 12710 3476 12716 3528
rect 12768 3476 12774 3528
rect 12989 3519 13047 3525
rect 12989 3485 13001 3519
rect 13035 3516 13047 3519
rect 13446 3516 13452 3528
rect 13035 3488 13452 3516
rect 13035 3485 13047 3488
rect 12989 3479 13047 3485
rect 13446 3476 13452 3488
rect 13504 3476 13510 3528
rect 13630 3476 13636 3528
rect 13688 3516 13694 3528
rect 13688 3488 15976 3516
rect 13688 3476 13694 3488
rect 9048 3420 9628 3448
rect 9858 3408 9864 3460
rect 9916 3448 9922 3460
rect 9916 3420 10640 3448
rect 9916 3408 9922 3420
rect 8018 3380 8024 3392
rect 7852 3352 8024 3380
rect 7745 3343 7803 3349
rect 8018 3340 8024 3352
rect 8076 3340 8082 3392
rect 8113 3383 8171 3389
rect 8113 3349 8125 3383
rect 8159 3380 8171 3383
rect 8202 3380 8208 3392
rect 8159 3352 8208 3380
rect 8159 3349 8171 3352
rect 8113 3343 8171 3349
rect 8202 3340 8208 3352
rect 8260 3340 8266 3392
rect 8389 3383 8447 3389
rect 8389 3349 8401 3383
rect 8435 3380 8447 3383
rect 8846 3380 8852 3392
rect 8435 3352 8852 3380
rect 8435 3349 8447 3352
rect 8389 3343 8447 3349
rect 8846 3340 8852 3352
rect 8904 3340 8910 3392
rect 10612 3380 10640 3420
rect 10870 3408 10876 3460
rect 10928 3448 10934 3460
rect 10928 3420 14596 3448
rect 10928 3408 10934 3420
rect 12066 3380 12072 3392
rect 10612 3352 12072 3380
rect 12066 3340 12072 3352
rect 12124 3340 12130 3392
rect 12437 3383 12495 3389
rect 12437 3349 12449 3383
rect 12483 3380 12495 3383
rect 12526 3380 12532 3392
rect 12483 3352 12532 3380
rect 12483 3349 12495 3352
rect 12437 3343 12495 3349
rect 12526 3340 12532 3352
rect 12584 3340 12590 3392
rect 12618 3340 12624 3392
rect 12676 3380 12682 3392
rect 13354 3380 13360 3392
rect 12676 3352 13360 3380
rect 12676 3340 12682 3352
rect 13354 3340 13360 3352
rect 13412 3340 13418 3392
rect 14568 3380 14596 3420
rect 15378 3408 15384 3460
rect 15436 3408 15442 3460
rect 15948 3448 15976 3488
rect 16022 3476 16028 3528
rect 16080 3476 16086 3528
rect 16132 3448 16160 3556
rect 16390 3476 16396 3528
rect 16448 3476 16454 3528
rect 16485 3519 16543 3525
rect 16485 3485 16497 3519
rect 16531 3485 16543 3519
rect 16485 3479 16543 3485
rect 15948 3420 16160 3448
rect 16298 3408 16304 3460
rect 16356 3448 16362 3460
rect 16500 3448 16528 3479
rect 16574 3476 16580 3528
rect 16632 3516 16638 3528
rect 16669 3519 16727 3525
rect 16669 3516 16681 3519
rect 16632 3488 16681 3516
rect 16632 3476 16638 3488
rect 16669 3485 16681 3488
rect 16715 3485 16727 3519
rect 16669 3479 16727 3485
rect 16850 3476 16856 3528
rect 16908 3476 16914 3528
rect 17052 3525 17080 3556
rect 17236 3525 17264 3624
rect 17402 3544 17408 3596
rect 17460 3544 17466 3596
rect 18046 3584 18052 3596
rect 17696 3556 18052 3584
rect 17037 3519 17095 3525
rect 17037 3485 17049 3519
rect 17083 3485 17095 3519
rect 17037 3479 17095 3485
rect 17221 3519 17279 3525
rect 17221 3485 17233 3519
rect 17267 3485 17279 3519
rect 17221 3479 17279 3485
rect 17310 3476 17316 3528
rect 17368 3476 17374 3528
rect 17494 3476 17500 3528
rect 17552 3516 17558 3528
rect 17696 3525 17724 3556
rect 18046 3544 18052 3556
rect 18104 3544 18110 3596
rect 17589 3519 17647 3525
rect 17589 3516 17601 3519
rect 17552 3488 17601 3516
rect 17552 3476 17558 3488
rect 17589 3485 17601 3488
rect 17635 3485 17647 3519
rect 17589 3479 17647 3485
rect 17681 3519 17739 3525
rect 17681 3485 17693 3519
rect 17727 3485 17739 3519
rect 17681 3479 17739 3485
rect 17954 3476 17960 3528
rect 18012 3476 18018 3528
rect 18138 3476 18144 3528
rect 18196 3476 18202 3528
rect 16356 3420 16528 3448
rect 16356 3408 16362 3420
rect 16761 3383 16819 3389
rect 16761 3380 16773 3383
rect 14568 3352 16773 3380
rect 16761 3349 16773 3352
rect 16807 3349 16819 3383
rect 16761 3343 16819 3349
rect 1104 3290 18860 3312
rect 1104 3238 2610 3290
rect 2662 3238 2674 3290
rect 2726 3238 2738 3290
rect 2790 3238 2802 3290
rect 2854 3238 2866 3290
rect 2918 3238 7610 3290
rect 7662 3238 7674 3290
rect 7726 3238 7738 3290
rect 7790 3238 7802 3290
rect 7854 3238 7866 3290
rect 7918 3238 12610 3290
rect 12662 3238 12674 3290
rect 12726 3238 12738 3290
rect 12790 3238 12802 3290
rect 12854 3238 12866 3290
rect 12918 3238 17610 3290
rect 17662 3238 17674 3290
rect 17726 3238 17738 3290
rect 17790 3238 17802 3290
rect 17854 3238 17866 3290
rect 17918 3238 18860 3290
rect 1104 3216 18860 3238
rect 3421 3179 3479 3185
rect 3421 3145 3433 3179
rect 3467 3176 3479 3179
rect 3694 3176 3700 3188
rect 3467 3148 3700 3176
rect 3467 3145 3479 3148
rect 3421 3139 3479 3145
rect 3694 3136 3700 3148
rect 3752 3136 3758 3188
rect 6730 3136 6736 3188
rect 6788 3176 6794 3188
rect 7466 3176 7472 3188
rect 6788 3148 7472 3176
rect 6788 3136 6794 3148
rect 7466 3136 7472 3148
rect 7524 3136 7530 3188
rect 8938 3136 8944 3188
rect 8996 3136 9002 3188
rect 10410 3176 10416 3188
rect 9508 3148 10416 3176
rect 1765 3111 1823 3117
rect 1765 3077 1777 3111
rect 1811 3108 1823 3111
rect 5166 3108 5172 3120
rect 1811 3080 5172 3108
rect 1811 3077 1823 3080
rect 1765 3071 1823 3077
rect 5166 3068 5172 3080
rect 5224 3068 5230 3120
rect 5353 3111 5411 3117
rect 5353 3077 5365 3111
rect 5399 3108 5411 3111
rect 5442 3108 5448 3120
rect 5399 3080 5448 3108
rect 5399 3077 5411 3080
rect 5353 3071 5411 3077
rect 5442 3068 5448 3080
rect 5500 3068 5506 3120
rect 7650 3108 7656 3120
rect 6288 3080 7656 3108
rect 2406 3000 2412 3052
rect 2464 3000 2470 3052
rect 2774 3000 2780 3052
rect 2832 3000 2838 3052
rect 2958 3000 2964 3052
rect 3016 3000 3022 3052
rect 3053 3043 3111 3049
rect 3053 3009 3065 3043
rect 3099 3040 3111 3043
rect 3326 3040 3332 3052
rect 3099 3012 3332 3040
rect 3099 3009 3111 3012
rect 3053 3003 3111 3009
rect 3326 3000 3332 3012
rect 3384 3000 3390 3052
rect 3510 3000 3516 3052
rect 3568 3000 3574 3052
rect 5718 3040 5724 3052
rect 3804 3012 5724 3040
rect 2225 2975 2283 2981
rect 2225 2941 2237 2975
rect 2271 2972 2283 2975
rect 2498 2972 2504 2984
rect 2271 2944 2504 2972
rect 2271 2941 2283 2944
rect 2225 2935 2283 2941
rect 2498 2932 2504 2944
rect 2556 2932 2562 2984
rect 2608 2944 3096 2972
rect 1581 2907 1639 2913
rect 1581 2873 1593 2907
rect 1627 2904 1639 2907
rect 2608 2904 2636 2944
rect 1627 2876 2636 2904
rect 2685 2907 2743 2913
rect 1627 2873 1639 2876
rect 1581 2867 1639 2873
rect 2685 2873 2697 2907
rect 2731 2873 2743 2907
rect 3068 2904 3096 2944
rect 3142 2932 3148 2984
rect 3200 2932 3206 2984
rect 3234 2932 3240 2984
rect 3292 2932 3298 2984
rect 3804 2904 3832 3012
rect 5718 3000 5724 3012
rect 5776 3000 5782 3052
rect 4246 2932 4252 2984
rect 4304 2972 4310 2984
rect 6288 2972 6316 3080
rect 7650 3068 7656 3080
rect 7708 3068 7714 3120
rect 6365 3043 6423 3049
rect 6365 3009 6377 3043
rect 6411 3009 6423 3043
rect 6365 3003 6423 3009
rect 4304 2944 6316 2972
rect 6380 2972 6408 3003
rect 6546 3000 6552 3052
rect 6604 3000 6610 3052
rect 6638 3000 6644 3052
rect 6696 3040 6702 3052
rect 6825 3043 6883 3049
rect 6825 3040 6837 3043
rect 6696 3012 6837 3040
rect 6696 3000 6702 3012
rect 6825 3009 6837 3012
rect 6871 3009 6883 3043
rect 8113 3043 8171 3049
rect 8113 3040 8125 3043
rect 6825 3003 6883 3009
rect 6932 3012 8125 3040
rect 6454 2972 6460 2984
rect 6380 2944 6460 2972
rect 4304 2932 4310 2944
rect 6454 2932 6460 2944
rect 6512 2932 6518 2984
rect 6932 2972 6960 3012
rect 8113 3009 8125 3012
rect 8159 3009 8171 3043
rect 8113 3003 8171 3009
rect 8294 3000 8300 3052
rect 8352 3000 8358 3052
rect 8386 3022 8392 3074
rect 8444 3022 8450 3074
rect 9122 3068 9128 3120
rect 9180 3108 9186 3120
rect 9180 3080 9444 3108
rect 9180 3068 9186 3080
rect 8481 3043 8539 3049
rect 8481 3009 8493 3043
rect 8527 3040 8539 3043
rect 8757 3043 8815 3049
rect 8527 3012 8708 3040
rect 8527 3009 8539 3012
rect 8481 3003 8539 3009
rect 6564 2944 6960 2972
rect 3068 2876 3832 2904
rect 2685 2867 2743 2873
rect 2700 2836 2728 2867
rect 3878 2864 3884 2916
rect 3936 2864 3942 2916
rect 5074 2864 5080 2916
rect 5132 2904 5138 2916
rect 6564 2904 6592 2944
rect 7926 2932 7932 2984
rect 7984 2932 7990 2984
rect 8570 2932 8576 2984
rect 8628 2932 8634 2984
rect 8680 2972 8708 3012
rect 8757 3009 8769 3043
rect 8803 3040 8815 3043
rect 8803 3012 9260 3040
rect 8803 3009 8815 3012
rect 8757 3003 8815 3009
rect 8846 2972 8852 2984
rect 8680 2944 8852 2972
rect 8846 2932 8852 2944
rect 8904 2932 8910 2984
rect 9232 2972 9260 3012
rect 9306 3000 9312 3052
rect 9364 3000 9370 3052
rect 9416 3049 9444 3080
rect 9401 3043 9459 3049
rect 9401 3009 9413 3043
rect 9447 3009 9459 3043
rect 9401 3003 9459 3009
rect 9508 2972 9536 3148
rect 10410 3136 10416 3148
rect 10468 3136 10474 3188
rect 11698 3185 11704 3188
rect 11685 3179 11704 3185
rect 11685 3145 11697 3179
rect 11756 3176 11762 3188
rect 14090 3176 14096 3188
rect 11756 3148 14096 3176
rect 11685 3139 11704 3145
rect 11698 3136 11704 3139
rect 11756 3136 11762 3148
rect 14090 3136 14096 3148
rect 14148 3136 14154 3188
rect 14458 3136 14464 3188
rect 14516 3176 14522 3188
rect 17402 3176 17408 3188
rect 14516 3148 17408 3176
rect 14516 3136 14522 3148
rect 17402 3136 17408 3148
rect 17460 3136 17466 3188
rect 9950 3108 9956 3120
rect 9600 3080 9956 3108
rect 9600 3052 9628 3080
rect 9950 3068 9956 3080
rect 10008 3068 10014 3120
rect 11054 3068 11060 3120
rect 11112 3108 11118 3120
rect 11333 3111 11391 3117
rect 11333 3108 11345 3111
rect 11112 3080 11345 3108
rect 11112 3068 11118 3080
rect 11333 3077 11345 3080
rect 11379 3077 11391 3111
rect 11333 3071 11391 3077
rect 11882 3068 11888 3120
rect 11940 3068 11946 3120
rect 12161 3111 12219 3117
rect 12161 3108 12173 3111
rect 11992 3080 12173 3108
rect 9582 3000 9588 3052
rect 9640 3000 9646 3052
rect 9769 3043 9827 3049
rect 9769 3009 9781 3043
rect 9815 3040 9827 3043
rect 10778 3040 10784 3052
rect 9815 3012 10784 3040
rect 9815 3009 9827 3012
rect 9769 3003 9827 3009
rect 10778 3000 10784 3012
rect 10836 3000 10842 3052
rect 10962 3000 10968 3052
rect 11020 3040 11026 3052
rect 11149 3043 11207 3049
rect 11149 3040 11161 3043
rect 11020 3012 11161 3040
rect 11020 3000 11026 3012
rect 11149 3009 11161 3012
rect 11195 3009 11207 3043
rect 11149 3003 11207 3009
rect 11606 3000 11612 3052
rect 11664 3040 11670 3052
rect 11992 3040 12020 3080
rect 12161 3077 12173 3080
rect 12207 3077 12219 3111
rect 12161 3071 12219 3077
rect 16206 3068 16212 3120
rect 16264 3108 16270 3120
rect 16264 3080 17448 3108
rect 16264 3068 16270 3080
rect 11664 3012 12020 3040
rect 11664 3000 11670 3012
rect 12066 3000 12072 3052
rect 12124 3000 12130 3052
rect 12253 3043 12311 3049
rect 12253 3009 12265 3043
rect 12299 3009 12311 3043
rect 12253 3003 12311 3009
rect 9232 2944 9536 2972
rect 11238 2932 11244 2984
rect 11296 2972 11302 2984
rect 12268 2972 12296 3003
rect 12434 3000 12440 3052
rect 12492 3040 12498 3052
rect 12492 3012 12848 3040
rect 12492 3000 12498 3012
rect 11296 2944 12296 2972
rect 11296 2932 11302 2944
rect 12710 2932 12716 2984
rect 12768 2932 12774 2984
rect 12820 2972 12848 3012
rect 13078 3000 13084 3052
rect 13136 3040 13142 3052
rect 13630 3040 13636 3052
rect 13136 3012 13636 3040
rect 13136 3000 13142 3012
rect 13630 3000 13636 3012
rect 13688 3000 13694 3052
rect 15838 3000 15844 3052
rect 15896 3040 15902 3052
rect 16482 3040 16488 3052
rect 15896 3012 16488 3040
rect 15896 3000 15902 3012
rect 16482 3000 16488 3012
rect 16540 3040 16546 3052
rect 17420 3049 17448 3080
rect 17221 3043 17279 3049
rect 17221 3040 17233 3043
rect 16540 3012 17233 3040
rect 16540 3000 16546 3012
rect 17221 3009 17233 3012
rect 17267 3009 17279 3043
rect 17221 3003 17279 3009
rect 17405 3043 17463 3049
rect 17405 3009 17417 3043
rect 17451 3009 17463 3043
rect 17405 3003 17463 3009
rect 13265 2975 13323 2981
rect 13265 2972 13277 2975
rect 12820 2944 13277 2972
rect 13265 2941 13277 2944
rect 13311 2941 13323 2975
rect 13265 2935 13323 2941
rect 16942 2932 16948 2984
rect 17000 2972 17006 2984
rect 17310 2972 17316 2984
rect 17000 2944 17316 2972
rect 17000 2932 17006 2944
rect 17310 2932 17316 2944
rect 17368 2932 17374 2984
rect 5132 2876 6592 2904
rect 5132 2864 5138 2876
rect 6638 2864 6644 2916
rect 6696 2864 6702 2916
rect 6730 2864 6736 2916
rect 6788 2864 6794 2916
rect 6840 2876 7972 2904
rect 2958 2836 2964 2848
rect 2700 2808 2964 2836
rect 2958 2796 2964 2808
rect 3016 2796 3022 2848
rect 3970 2796 3976 2848
rect 4028 2796 4034 2848
rect 4890 2796 4896 2848
rect 4948 2836 4954 2848
rect 5261 2839 5319 2845
rect 5261 2836 5273 2839
rect 4948 2808 5273 2836
rect 4948 2796 4954 2808
rect 5261 2805 5273 2808
rect 5307 2836 5319 2839
rect 6546 2836 6552 2848
rect 5307 2808 6552 2836
rect 5307 2805 5319 2808
rect 5261 2799 5319 2805
rect 6546 2796 6552 2808
rect 6604 2836 6610 2848
rect 6840 2836 6868 2876
rect 6604 2808 6868 2836
rect 7009 2839 7067 2845
rect 6604 2796 6610 2808
rect 7009 2805 7021 2839
rect 7055 2836 7067 2839
rect 7834 2836 7840 2848
rect 7055 2808 7840 2836
rect 7055 2805 7067 2808
rect 7009 2799 7067 2805
rect 7834 2796 7840 2808
rect 7892 2796 7898 2848
rect 7944 2836 7972 2876
rect 8202 2864 8208 2916
rect 8260 2904 8266 2916
rect 8260 2876 11744 2904
rect 8260 2864 8266 2876
rect 10594 2836 10600 2848
rect 7944 2808 10600 2836
rect 10594 2796 10600 2808
rect 10652 2836 10658 2848
rect 10778 2836 10784 2848
rect 10652 2808 10784 2836
rect 10652 2796 10658 2808
rect 10778 2796 10784 2808
rect 10836 2796 10842 2848
rect 11057 2839 11115 2845
rect 11057 2805 11069 2839
rect 11103 2836 11115 2839
rect 11330 2836 11336 2848
rect 11103 2808 11336 2836
rect 11103 2805 11115 2808
rect 11057 2799 11115 2805
rect 11330 2796 11336 2808
rect 11388 2796 11394 2848
rect 11517 2839 11575 2845
rect 11517 2805 11529 2839
rect 11563 2836 11575 2839
rect 11606 2836 11612 2848
rect 11563 2808 11612 2836
rect 11563 2805 11575 2808
rect 11517 2799 11575 2805
rect 11606 2796 11612 2808
rect 11664 2796 11670 2848
rect 11716 2845 11744 2876
rect 12342 2864 12348 2916
rect 12400 2904 12406 2916
rect 12805 2907 12863 2913
rect 12805 2904 12817 2907
rect 12400 2876 12817 2904
rect 12400 2864 12406 2876
rect 12805 2873 12817 2876
rect 12851 2873 12863 2907
rect 12805 2867 12863 2873
rect 13354 2864 13360 2916
rect 13412 2904 13418 2916
rect 18046 2904 18052 2916
rect 13412 2876 18052 2904
rect 13412 2864 13418 2876
rect 18046 2864 18052 2876
rect 18104 2864 18110 2916
rect 11701 2839 11759 2845
rect 11701 2805 11713 2839
rect 11747 2836 11759 2839
rect 14182 2836 14188 2848
rect 11747 2808 14188 2836
rect 11747 2805 11759 2808
rect 11701 2799 11759 2805
rect 14182 2796 14188 2808
rect 14240 2796 14246 2848
rect 16850 2796 16856 2848
rect 16908 2836 16914 2848
rect 17313 2839 17371 2845
rect 17313 2836 17325 2839
rect 16908 2808 17325 2836
rect 16908 2796 16914 2808
rect 17313 2805 17325 2808
rect 17359 2805 17371 2839
rect 17313 2799 17371 2805
rect 1104 2746 18860 2768
rect 1104 2694 1950 2746
rect 2002 2694 2014 2746
rect 2066 2694 2078 2746
rect 2130 2694 2142 2746
rect 2194 2694 2206 2746
rect 2258 2694 6950 2746
rect 7002 2694 7014 2746
rect 7066 2694 7078 2746
rect 7130 2694 7142 2746
rect 7194 2694 7206 2746
rect 7258 2694 11950 2746
rect 12002 2694 12014 2746
rect 12066 2694 12078 2746
rect 12130 2694 12142 2746
rect 12194 2694 12206 2746
rect 12258 2694 16950 2746
rect 17002 2694 17014 2746
rect 17066 2694 17078 2746
rect 17130 2694 17142 2746
rect 17194 2694 17206 2746
rect 17258 2694 18860 2746
rect 1104 2672 18860 2694
rect 1670 2592 1676 2644
rect 1728 2632 1734 2644
rect 2317 2635 2375 2641
rect 2317 2632 2329 2635
rect 1728 2604 2329 2632
rect 1728 2592 1734 2604
rect 2317 2601 2329 2604
rect 2363 2601 2375 2635
rect 2317 2595 2375 2601
rect 2777 2635 2835 2641
rect 2777 2601 2789 2635
rect 2823 2632 2835 2635
rect 3418 2632 3424 2644
rect 2823 2604 3424 2632
rect 2823 2601 2835 2604
rect 2777 2595 2835 2601
rect 3418 2592 3424 2604
rect 3476 2592 3482 2644
rect 3786 2592 3792 2644
rect 3844 2632 3850 2644
rect 3973 2635 4031 2641
rect 3973 2632 3985 2635
rect 3844 2604 3985 2632
rect 3844 2592 3850 2604
rect 3973 2601 3985 2604
rect 4019 2601 4031 2635
rect 3973 2595 4031 2601
rect 5442 2592 5448 2644
rect 5500 2632 5506 2644
rect 6641 2635 6699 2641
rect 6641 2632 6653 2635
rect 5500 2604 6653 2632
rect 5500 2592 5506 2604
rect 6641 2601 6653 2604
rect 6687 2601 6699 2635
rect 6641 2595 6699 2601
rect 9030 2592 9036 2644
rect 9088 2592 9094 2644
rect 9214 2592 9220 2644
rect 9272 2632 9278 2644
rect 13354 2632 13360 2644
rect 9272 2604 10364 2632
rect 9272 2592 9278 2604
rect 1964 2536 6224 2564
rect 474 2456 480 2508
rect 532 2496 538 2508
rect 1397 2499 1455 2505
rect 1397 2496 1409 2499
rect 532 2468 1409 2496
rect 532 2456 538 2468
rect 1228 2292 1256 2468
rect 1397 2465 1409 2468
rect 1443 2465 1455 2499
rect 1397 2459 1455 2465
rect 1302 2388 1308 2440
rect 1360 2428 1366 2440
rect 1360 2400 1532 2428
rect 1360 2388 1366 2400
rect 1504 2360 1532 2400
rect 1670 2388 1676 2440
rect 1728 2428 1734 2440
rect 1854 2428 1860 2440
rect 1728 2400 1860 2428
rect 1728 2388 1734 2400
rect 1854 2388 1860 2400
rect 1912 2388 1918 2440
rect 1964 2437 1992 2536
rect 2501 2499 2559 2505
rect 2501 2465 2513 2499
rect 2547 2496 2559 2499
rect 4982 2496 4988 2508
rect 2547 2468 4988 2496
rect 2547 2465 2559 2468
rect 2501 2459 2559 2465
rect 4982 2456 4988 2468
rect 5040 2456 5046 2508
rect 6196 2496 6224 2536
rect 6546 2524 6552 2576
rect 6604 2564 6610 2576
rect 9306 2564 9312 2576
rect 6604 2536 9312 2564
rect 6604 2524 6610 2536
rect 9306 2524 9312 2536
rect 9364 2524 9370 2576
rect 10336 2564 10364 2604
rect 10520 2604 13360 2632
rect 10520 2564 10548 2604
rect 13354 2592 13360 2604
rect 13412 2592 13418 2644
rect 10336 2536 10548 2564
rect 11422 2524 11428 2576
rect 11480 2564 11486 2576
rect 12805 2567 12863 2573
rect 12805 2564 12817 2567
rect 11480 2536 12817 2564
rect 11480 2524 11486 2536
rect 12805 2533 12817 2536
rect 12851 2533 12863 2567
rect 12805 2527 12863 2533
rect 6730 2496 6736 2508
rect 6196 2468 6736 2496
rect 6730 2456 6736 2468
rect 6788 2456 6794 2508
rect 7466 2456 7472 2508
rect 7524 2496 7530 2508
rect 8113 2499 8171 2505
rect 8113 2496 8125 2499
rect 7524 2468 8125 2496
rect 7524 2456 7530 2468
rect 8113 2465 8125 2468
rect 8159 2465 8171 2499
rect 8478 2496 8484 2508
rect 8113 2459 8171 2465
rect 8220 2468 8484 2496
rect 1949 2431 2007 2437
rect 1949 2397 1961 2431
rect 1995 2397 2007 2431
rect 1949 2391 2007 2397
rect 2038 2388 2044 2440
rect 2096 2388 2102 2440
rect 2225 2431 2283 2437
rect 2225 2397 2237 2431
rect 2271 2397 2283 2431
rect 2225 2391 2283 2397
rect 2240 2360 2268 2391
rect 2406 2388 2412 2440
rect 2464 2428 2470 2440
rect 2593 2431 2651 2437
rect 2593 2428 2605 2431
rect 2464 2400 2605 2428
rect 2464 2388 2470 2400
rect 2593 2397 2605 2400
rect 2639 2397 2651 2431
rect 4246 2428 4252 2440
rect 2593 2391 2651 2397
rect 3252 2400 4252 2428
rect 3252 2360 3280 2400
rect 4246 2388 4252 2400
rect 4304 2388 4310 2440
rect 6546 2388 6552 2440
rect 6604 2388 6610 2440
rect 7068 2431 7126 2437
rect 7068 2397 7080 2431
rect 7114 2428 7126 2431
rect 8220 2428 8248 2468
rect 8478 2456 8484 2468
rect 8536 2456 8542 2508
rect 8570 2456 8576 2508
rect 8628 2456 8634 2508
rect 8662 2456 8668 2508
rect 8720 2456 8726 2508
rect 9398 2456 9404 2508
rect 9456 2496 9462 2508
rect 9493 2499 9551 2505
rect 9493 2496 9505 2499
rect 9456 2468 9505 2496
rect 9456 2456 9462 2468
rect 9493 2465 9505 2468
rect 9539 2465 9551 2499
rect 9493 2459 9551 2465
rect 10413 2499 10471 2505
rect 10413 2465 10425 2499
rect 10459 2496 10471 2499
rect 11054 2496 11060 2508
rect 10459 2468 11060 2496
rect 10459 2465 10471 2468
rect 10413 2459 10471 2465
rect 11054 2456 11060 2468
rect 11112 2456 11118 2508
rect 12345 2499 12403 2505
rect 12345 2465 12357 2499
rect 12391 2496 12403 2499
rect 13814 2496 13820 2508
rect 12391 2468 13820 2496
rect 12391 2465 12403 2468
rect 12345 2459 12403 2465
rect 13814 2456 13820 2468
rect 13872 2456 13878 2508
rect 15286 2456 15292 2508
rect 15344 2496 15350 2508
rect 18506 2496 18512 2508
rect 15344 2468 18512 2496
rect 15344 2456 15350 2468
rect 18506 2456 18512 2468
rect 18564 2456 18570 2508
rect 7114 2400 8248 2428
rect 8297 2431 8355 2437
rect 7114 2397 7126 2400
rect 7068 2391 7126 2397
rect 8297 2397 8309 2431
rect 8343 2428 8355 2431
rect 8754 2428 8760 2440
rect 8343 2400 8760 2428
rect 8343 2397 8355 2400
rect 8297 2391 8355 2397
rect 8754 2388 8760 2400
rect 8812 2388 8818 2440
rect 9214 2388 9220 2440
rect 9272 2388 9278 2440
rect 9306 2388 9312 2440
rect 9364 2388 9370 2440
rect 9582 2388 9588 2440
rect 9640 2388 9646 2440
rect 10870 2428 10876 2440
rect 9692 2400 10876 2428
rect 1504 2332 2268 2360
rect 2424 2332 3280 2360
rect 2424 2292 2452 2332
rect 3326 2320 3332 2372
rect 3384 2360 3390 2372
rect 3881 2363 3939 2369
rect 3881 2360 3893 2363
rect 3384 2332 3893 2360
rect 3384 2320 3390 2332
rect 3881 2329 3893 2332
rect 3927 2329 3939 2363
rect 3881 2323 3939 2329
rect 8202 2320 8208 2372
rect 8260 2360 8266 2372
rect 9692 2360 9720 2400
rect 10870 2388 10876 2400
rect 10928 2388 10934 2440
rect 11146 2388 11152 2440
rect 11204 2388 11210 2440
rect 11330 2388 11336 2440
rect 11388 2388 11394 2440
rect 11606 2388 11612 2440
rect 11664 2388 11670 2440
rect 11698 2388 11704 2440
rect 11756 2428 11762 2440
rect 11793 2431 11851 2437
rect 11793 2428 11805 2431
rect 11756 2400 11805 2428
rect 11756 2388 11762 2400
rect 11793 2397 11805 2400
rect 11839 2397 11851 2431
rect 11793 2391 11851 2397
rect 11974 2388 11980 2440
rect 12032 2388 12038 2440
rect 12069 2431 12127 2437
rect 12069 2397 12081 2431
rect 12115 2428 12127 2431
rect 12434 2428 12440 2440
rect 12115 2400 12440 2428
rect 12115 2397 12127 2400
rect 12069 2391 12127 2397
rect 12434 2388 12440 2400
rect 12492 2388 12498 2440
rect 12621 2431 12679 2437
rect 12621 2397 12633 2431
rect 12667 2428 12679 2431
rect 12802 2428 12808 2440
rect 12667 2400 12808 2428
rect 12667 2397 12679 2400
rect 12621 2391 12679 2397
rect 12802 2388 12808 2400
rect 12860 2388 12866 2440
rect 12897 2431 12955 2437
rect 12897 2397 12909 2431
rect 12943 2428 12955 2431
rect 13722 2428 13728 2440
rect 12943 2400 13728 2428
rect 12943 2397 12955 2400
rect 12897 2391 12955 2397
rect 13722 2388 13728 2400
rect 13780 2388 13786 2440
rect 16574 2388 16580 2440
rect 16632 2428 16638 2440
rect 16669 2431 16727 2437
rect 16669 2428 16681 2431
rect 16632 2400 16681 2428
rect 16632 2388 16638 2400
rect 16669 2397 16681 2400
rect 16715 2397 16727 2431
rect 16669 2391 16727 2397
rect 16942 2388 16948 2440
rect 17000 2428 17006 2440
rect 17497 2431 17555 2437
rect 17497 2428 17509 2431
rect 17000 2400 17509 2428
rect 17000 2388 17006 2400
rect 17497 2397 17509 2400
rect 17543 2397 17555 2431
rect 17497 2391 17555 2397
rect 8260 2332 9720 2360
rect 8260 2320 8266 2332
rect 9950 2320 9956 2372
rect 10008 2360 10014 2372
rect 10137 2363 10195 2369
rect 10137 2360 10149 2363
rect 10008 2332 10149 2360
rect 10008 2320 10014 2332
rect 10137 2329 10149 2332
rect 10183 2329 10195 2363
rect 11624 2360 11652 2388
rect 15654 2360 15660 2372
rect 11624 2332 15660 2360
rect 10137 2323 10195 2329
rect 15654 2320 15660 2332
rect 15712 2320 15718 2372
rect 18322 2320 18328 2372
rect 18380 2320 18386 2372
rect 1228 2264 2452 2292
rect 2498 2252 2504 2304
rect 2556 2252 2562 2304
rect 4522 2252 4528 2304
rect 4580 2292 4586 2304
rect 7009 2295 7067 2301
rect 7009 2292 7021 2295
rect 4580 2264 7021 2292
rect 4580 2252 4586 2264
rect 7009 2261 7021 2264
rect 7055 2261 7067 2295
rect 7009 2255 7067 2261
rect 7190 2252 7196 2304
rect 7248 2252 7254 2304
rect 7650 2252 7656 2304
rect 7708 2292 7714 2304
rect 9122 2292 9128 2304
rect 7708 2264 9128 2292
rect 7708 2252 7714 2264
rect 9122 2252 9128 2264
rect 9180 2252 9186 2304
rect 11054 2252 11060 2304
rect 11112 2292 11118 2304
rect 11149 2295 11207 2301
rect 11149 2292 11161 2295
rect 11112 2264 11161 2292
rect 11112 2252 11118 2264
rect 11149 2261 11161 2264
rect 11195 2261 11207 2295
rect 11149 2255 11207 2261
rect 11606 2252 11612 2304
rect 11664 2252 11670 2304
rect 12434 2252 12440 2304
rect 12492 2292 12498 2304
rect 13262 2292 13268 2304
rect 12492 2264 13268 2292
rect 12492 2252 12498 2264
rect 13262 2252 13268 2264
rect 13320 2252 13326 2304
rect 16850 2252 16856 2304
rect 16908 2252 16914 2304
rect 1104 2202 18860 2224
rect 1104 2150 2610 2202
rect 2662 2150 2674 2202
rect 2726 2150 2738 2202
rect 2790 2150 2802 2202
rect 2854 2150 2866 2202
rect 2918 2150 7610 2202
rect 7662 2150 7674 2202
rect 7726 2150 7738 2202
rect 7790 2150 7802 2202
rect 7854 2150 7866 2202
rect 7918 2150 12610 2202
rect 12662 2150 12674 2202
rect 12726 2150 12738 2202
rect 12790 2150 12802 2202
rect 12854 2150 12866 2202
rect 12918 2150 17610 2202
rect 17662 2150 17674 2202
rect 17726 2150 17738 2202
rect 17790 2150 17802 2202
rect 17854 2150 17866 2202
rect 17918 2150 18860 2202
rect 1104 2128 18860 2150
rect 6730 2048 6736 2100
rect 6788 2088 6794 2100
rect 9398 2088 9404 2100
rect 6788 2060 9404 2088
rect 6788 2048 6794 2060
rect 9398 2048 9404 2060
rect 9456 2048 9462 2100
rect 10778 2048 10784 2100
rect 10836 2088 10842 2100
rect 13170 2088 13176 2100
rect 10836 2060 13176 2088
rect 10836 2048 10842 2060
rect 13170 2048 13176 2060
rect 13228 2048 13234 2100
rect 842 1980 848 2032
rect 900 2020 906 2032
rect 9214 2020 9220 2032
rect 900 1992 9220 2020
rect 900 1980 906 1992
rect 9214 1980 9220 1992
rect 9272 1980 9278 2032
rect 10962 1980 10968 2032
rect 11020 2020 11026 2032
rect 13538 2020 13544 2032
rect 11020 1992 13544 2020
rect 11020 1980 11026 1992
rect 13538 1980 13544 1992
rect 13596 2020 13602 2032
rect 16850 2020 16856 2032
rect 13596 1992 16856 2020
rect 13596 1980 13602 1992
rect 16850 1980 16856 1992
rect 16908 1980 16914 2032
rect 4062 1912 4068 1964
rect 4120 1952 4126 1964
rect 10686 1952 10692 1964
rect 4120 1924 10692 1952
rect 4120 1912 4126 1924
rect 10686 1912 10692 1924
rect 10744 1912 10750 1964
rect 9306 1844 9312 1896
rect 9364 1884 9370 1896
rect 17954 1884 17960 1896
rect 9364 1856 17960 1884
rect 9364 1844 9370 1856
rect 17954 1844 17960 1856
rect 18012 1844 18018 1896
rect 3050 1776 3056 1828
rect 3108 1816 3114 1828
rect 11514 1816 11520 1828
rect 3108 1788 11520 1816
rect 3108 1776 3114 1788
rect 11514 1776 11520 1788
rect 11572 1776 11578 1828
rect 7466 1708 7472 1760
rect 7524 1748 7530 1760
rect 11054 1748 11060 1760
rect 7524 1720 11060 1748
rect 7524 1708 7530 1720
rect 11054 1708 11060 1720
rect 11112 1708 11118 1760
rect 14918 1748 14924 1760
rect 12406 1720 14924 1748
rect 1670 1640 1676 1692
rect 1728 1680 1734 1692
rect 6454 1680 6460 1692
rect 1728 1652 6460 1680
rect 1728 1640 1734 1652
rect 6454 1640 6460 1652
rect 6512 1680 6518 1692
rect 12406 1680 12434 1720
rect 14918 1708 14924 1720
rect 14976 1708 14982 1760
rect 6512 1652 12434 1680
rect 6512 1640 6518 1652
rect 6270 1572 6276 1624
rect 6328 1612 6334 1624
rect 9766 1612 9772 1624
rect 6328 1584 9772 1612
rect 6328 1572 6334 1584
rect 9766 1572 9772 1584
rect 9824 1572 9830 1624
rect 8478 1504 8484 1556
rect 8536 1544 8542 1556
rect 17494 1544 17500 1556
rect 8536 1516 17500 1544
rect 8536 1504 8542 1516
rect 17494 1504 17500 1516
rect 17552 1504 17558 1556
rect 5718 1436 5724 1488
rect 5776 1476 5782 1488
rect 13078 1476 13084 1488
rect 5776 1448 13084 1476
rect 5776 1436 5782 1448
rect 13078 1436 13084 1448
rect 13136 1436 13142 1488
rect 2314 1300 2320 1352
rect 2372 1340 2378 1352
rect 6086 1340 6092 1352
rect 2372 1312 6092 1340
rect 2372 1300 2378 1312
rect 6086 1300 6092 1312
rect 6144 1300 6150 1352
rect 6178 1300 6184 1352
rect 6236 1340 6242 1352
rect 11146 1340 11152 1352
rect 6236 1312 11152 1340
rect 6236 1300 6242 1312
rect 11146 1300 11152 1312
rect 11204 1300 11210 1352
rect 4614 1232 4620 1284
rect 4672 1272 4678 1284
rect 11238 1272 11244 1284
rect 4672 1244 11244 1272
rect 4672 1232 4678 1244
rect 11238 1232 11244 1244
rect 11296 1232 11302 1284
rect 12986 1272 12992 1284
rect 11348 1244 12992 1272
rect 7282 1164 7288 1216
rect 7340 1204 7346 1216
rect 11348 1204 11376 1244
rect 12986 1232 12992 1244
rect 13044 1232 13050 1284
rect 16758 1204 16764 1216
rect 7340 1176 11376 1204
rect 12406 1176 16764 1204
rect 7340 1164 7346 1176
rect 6362 1096 6368 1148
rect 6420 1136 6426 1148
rect 12406 1136 12434 1176
rect 16758 1164 16764 1176
rect 16816 1164 16822 1216
rect 6420 1108 12434 1136
rect 6420 1096 6426 1108
rect 2958 1028 2964 1080
rect 3016 1068 3022 1080
rect 5810 1068 5816 1080
rect 3016 1040 5816 1068
rect 3016 1028 3022 1040
rect 5810 1028 5816 1040
rect 5868 1068 5874 1080
rect 16022 1068 16028 1080
rect 5868 1040 16028 1068
rect 5868 1028 5874 1040
rect 16022 1028 16028 1040
rect 16080 1028 16086 1080
rect 4154 960 4160 1012
rect 4212 1000 4218 1012
rect 11790 1000 11796 1012
rect 4212 972 11796 1000
rect 4212 960 4218 972
rect 11790 960 11796 972
rect 11848 960 11854 1012
rect 3142 892 3148 944
rect 3200 932 3206 944
rect 15378 932 15384 944
rect 3200 904 15384 932
rect 3200 892 3206 904
rect 15378 892 15384 904
rect 15436 892 15442 944
rect 5994 824 6000 876
rect 6052 864 6058 876
rect 15470 864 15476 876
rect 6052 836 15476 864
rect 6052 824 6058 836
rect 15470 824 15476 836
rect 15528 824 15534 876
rect 5166 756 5172 808
rect 5224 796 5230 808
rect 17310 796 17316 808
rect 5224 768 17316 796
rect 5224 756 5230 768
rect 17310 756 17316 768
rect 17368 756 17374 808
rect 5258 620 5264 672
rect 5316 660 5322 672
rect 12526 660 12532 672
rect 5316 632 12532 660
rect 5316 620 5322 632
rect 12526 620 12532 632
rect 12584 620 12590 672
rect 6638 552 6644 604
rect 6696 592 6702 604
rect 14274 592 14280 604
rect 6696 564 14280 592
rect 6696 552 6702 564
rect 14274 552 14280 564
rect 14332 552 14338 604
rect 3970 484 3976 536
rect 4028 524 4034 536
rect 14642 524 14648 536
rect 4028 496 14648 524
rect 4028 484 4034 496
rect 14642 484 14648 496
rect 14700 484 14706 536
<< via1 >>
rect 5816 18776 5868 18828
rect 11520 18776 11572 18828
rect 6092 18708 6144 18760
rect 14280 18708 14332 18760
rect 1584 18572 1636 18624
rect 10232 18572 10284 18624
rect 5632 18504 5684 18556
rect 15936 18504 15988 18556
rect 3332 18436 3384 18488
rect 14464 18436 14516 18488
rect 9680 18368 9732 18420
rect 11428 18368 11480 18420
rect 11520 18368 11572 18420
rect 16764 18368 16816 18420
rect 5264 18300 5316 18352
rect 14648 18300 14700 18352
rect 8576 18232 8628 18284
rect 14372 18232 14424 18284
rect 6736 18164 6788 18216
rect 11428 18164 11480 18216
rect 16304 18164 16356 18216
rect 13820 18096 13872 18148
rect 9036 18028 9088 18080
rect 15292 18028 15344 18080
rect 3608 17960 3660 18012
rect 10784 17960 10836 18012
rect 4436 17756 4488 17808
rect 9588 17756 9640 17808
rect 15936 17756 15988 17808
rect 19524 17756 19576 17808
rect 4804 17688 4856 17740
rect 9864 17688 9916 17740
rect 3976 17620 4028 17672
rect 16488 17620 16540 17672
rect 8208 17552 8260 17604
rect 15384 17552 15436 17604
rect 3516 17484 3568 17536
rect 9772 17484 9824 17536
rect 9864 17484 9916 17536
rect 16672 17484 16724 17536
rect 2610 17382 2662 17434
rect 2674 17382 2726 17434
rect 2738 17382 2790 17434
rect 2802 17382 2854 17434
rect 2866 17382 2918 17434
rect 7610 17382 7662 17434
rect 7674 17382 7726 17434
rect 7738 17382 7790 17434
rect 7802 17382 7854 17434
rect 7866 17382 7918 17434
rect 12610 17382 12662 17434
rect 12674 17382 12726 17434
rect 12738 17382 12790 17434
rect 12802 17382 12854 17434
rect 12866 17382 12918 17434
rect 17610 17382 17662 17434
rect 17674 17382 17726 17434
rect 17738 17382 17790 17434
rect 17802 17382 17854 17434
rect 17866 17382 17918 17434
rect 940 17280 992 17332
rect 9496 17280 9548 17332
rect 15660 17280 15712 17332
rect 17500 17280 17552 17332
rect 2964 17212 3016 17264
rect 3700 17212 3752 17264
rect 3056 17144 3108 17196
rect 5448 17187 5500 17196
rect 5448 17153 5457 17187
rect 5457 17153 5491 17187
rect 5491 17153 5500 17187
rect 5448 17144 5500 17153
rect 6184 17212 6236 17264
rect 8668 17212 8720 17264
rect 9772 17255 9824 17264
rect 9772 17221 9781 17255
rect 9781 17221 9815 17255
rect 9815 17221 9824 17255
rect 9772 17212 9824 17221
rect 7380 17144 7432 17196
rect 13176 17212 13228 17264
rect 5356 17119 5408 17128
rect 5356 17085 5365 17119
rect 5365 17085 5399 17119
rect 5399 17085 5408 17119
rect 5356 17076 5408 17085
rect 11152 17144 11204 17196
rect 9588 17076 9640 17128
rect 10508 17076 10560 17128
rect 13636 17144 13688 17196
rect 16120 17144 16172 17196
rect 17316 17187 17368 17196
rect 17316 17153 17325 17187
rect 17325 17153 17359 17187
rect 17359 17153 17368 17187
rect 17316 17144 17368 17153
rect 18604 17144 18656 17196
rect 10416 17008 10468 17060
rect 11980 17076 12032 17128
rect 16028 17119 16080 17128
rect 16028 17085 16037 17119
rect 16037 17085 16071 17119
rect 16071 17085 16080 17119
rect 16028 17076 16080 17085
rect 18144 17076 18196 17128
rect 1768 16983 1820 16992
rect 1768 16949 1777 16983
rect 1777 16949 1811 16983
rect 1811 16949 1820 16983
rect 1768 16940 1820 16949
rect 2412 16940 2464 16992
rect 4896 16940 4948 16992
rect 6276 16940 6328 16992
rect 8760 16940 8812 16992
rect 17316 17008 17368 17060
rect 11336 16940 11388 16992
rect 12992 16940 13044 16992
rect 1950 16838 2002 16890
rect 2014 16838 2066 16890
rect 2078 16838 2130 16890
rect 2142 16838 2194 16890
rect 2206 16838 2258 16890
rect 6950 16838 7002 16890
rect 7014 16838 7066 16890
rect 7078 16838 7130 16890
rect 7142 16838 7194 16890
rect 7206 16838 7258 16890
rect 11950 16838 12002 16890
rect 12014 16838 12066 16890
rect 12078 16838 12130 16890
rect 12142 16838 12194 16890
rect 12206 16838 12258 16890
rect 16950 16838 17002 16890
rect 17014 16838 17066 16890
rect 17078 16838 17130 16890
rect 17142 16838 17194 16890
rect 17206 16838 17258 16890
rect 8116 16736 8168 16788
rect 13544 16736 13596 16788
rect 13728 16736 13780 16788
rect 4988 16668 5040 16720
rect 10508 16668 10560 16720
rect 10692 16711 10744 16720
rect 10692 16677 10701 16711
rect 10701 16677 10735 16711
rect 10735 16677 10744 16711
rect 10692 16668 10744 16677
rect 10784 16668 10836 16720
rect 1860 16600 1912 16652
rect 5448 16600 5500 16652
rect 8576 16600 8628 16652
rect 8852 16600 8904 16652
rect 12440 16600 12492 16652
rect 15200 16643 15252 16652
rect 15200 16609 15209 16643
rect 15209 16609 15243 16643
rect 15243 16609 15252 16643
rect 15200 16600 15252 16609
rect 15568 16736 15620 16788
rect 16212 16668 16264 16720
rect 1216 16532 1268 16584
rect 10416 16575 10468 16584
rect 10416 16541 10425 16575
rect 10425 16541 10459 16575
rect 10459 16541 10468 16575
rect 10416 16532 10468 16541
rect 10600 16532 10652 16584
rect 11612 16532 11664 16584
rect 16120 16532 16172 16584
rect 17040 16575 17092 16584
rect 17040 16541 17049 16575
rect 17049 16541 17083 16575
rect 17083 16541 17092 16575
rect 17040 16532 17092 16541
rect 17132 16575 17184 16584
rect 17132 16541 17141 16575
rect 17141 16541 17175 16575
rect 17175 16541 17184 16575
rect 17132 16532 17184 16541
rect 1492 16507 1544 16516
rect 1492 16473 1501 16507
rect 1501 16473 1535 16507
rect 1535 16473 1544 16507
rect 1492 16464 1544 16473
rect 3148 16464 3200 16516
rect 11336 16464 11388 16516
rect 11520 16464 11572 16516
rect 13452 16464 13504 16516
rect 14188 16464 14240 16516
rect 16396 16507 16448 16516
rect 16396 16473 16405 16507
rect 16405 16473 16439 16507
rect 16439 16473 16448 16507
rect 16396 16464 16448 16473
rect 10508 16439 10560 16448
rect 10508 16405 10517 16439
rect 10517 16405 10551 16439
rect 10551 16405 10560 16439
rect 10508 16396 10560 16405
rect 10876 16396 10928 16448
rect 17960 16464 18012 16516
rect 16764 16396 16816 16448
rect 18420 16439 18472 16448
rect 18420 16405 18429 16439
rect 18429 16405 18463 16439
rect 18463 16405 18472 16439
rect 18420 16396 18472 16405
rect 2610 16294 2662 16346
rect 2674 16294 2726 16346
rect 2738 16294 2790 16346
rect 2802 16294 2854 16346
rect 2866 16294 2918 16346
rect 7610 16294 7662 16346
rect 7674 16294 7726 16346
rect 7738 16294 7790 16346
rect 7802 16294 7854 16346
rect 7866 16294 7918 16346
rect 12610 16294 12662 16346
rect 12674 16294 12726 16346
rect 12738 16294 12790 16346
rect 12802 16294 12854 16346
rect 12866 16294 12918 16346
rect 17610 16294 17662 16346
rect 17674 16294 17726 16346
rect 17738 16294 17790 16346
rect 17802 16294 17854 16346
rect 17866 16294 17918 16346
rect 4620 16192 4672 16244
rect 5172 16192 5224 16244
rect 12992 16192 13044 16244
rect 17132 16192 17184 16244
rect 2780 15988 2832 16040
rect 848 15920 900 15972
rect 7380 16124 7432 16176
rect 9128 16124 9180 16176
rect 3056 16099 3108 16108
rect 3056 16065 3065 16099
rect 3065 16065 3099 16099
rect 3099 16065 3108 16099
rect 3056 16056 3108 16065
rect 6552 16099 6604 16108
rect 6552 16065 6561 16099
rect 6561 16065 6595 16099
rect 6595 16065 6604 16099
rect 6552 16056 6604 16065
rect 6644 16099 6696 16108
rect 6644 16065 6653 16099
rect 6653 16065 6687 16099
rect 6687 16065 6696 16099
rect 6644 16056 6696 16065
rect 7012 16099 7064 16108
rect 7012 16065 7021 16099
rect 7021 16065 7055 16099
rect 7055 16065 7064 16099
rect 7012 16056 7064 16065
rect 7840 16056 7892 16108
rect 8208 16056 8260 16108
rect 9220 16056 9272 16108
rect 12532 16124 12584 16176
rect 13544 16124 13596 16176
rect 18236 16124 18288 16176
rect 12624 16099 12676 16108
rect 6460 15988 6512 16040
rect 7748 15988 7800 16040
rect 10416 15988 10468 16040
rect 10876 15988 10928 16040
rect 11612 15988 11664 16040
rect 12624 16065 12633 16099
rect 12633 16065 12667 16099
rect 12667 16065 12676 16099
rect 12624 16056 12676 16065
rect 16580 16056 16632 16108
rect 17500 15988 17552 16040
rect 4160 15920 4212 15972
rect 10048 15920 10100 15972
rect 10692 15920 10744 15972
rect 12532 15920 12584 15972
rect 7380 15852 7432 15904
rect 8024 15852 8076 15904
rect 10324 15852 10376 15904
rect 11612 15852 11664 15904
rect 18788 15852 18840 15904
rect 1950 15750 2002 15802
rect 2014 15750 2066 15802
rect 2078 15750 2130 15802
rect 2142 15750 2194 15802
rect 2206 15750 2258 15802
rect 6950 15750 7002 15802
rect 7014 15750 7066 15802
rect 7078 15750 7130 15802
rect 7142 15750 7194 15802
rect 7206 15750 7258 15802
rect 11950 15750 12002 15802
rect 12014 15750 12066 15802
rect 12078 15750 12130 15802
rect 12142 15750 12194 15802
rect 12206 15750 12258 15802
rect 16950 15750 17002 15802
rect 17014 15750 17066 15802
rect 17078 15750 17130 15802
rect 17142 15750 17194 15802
rect 17206 15750 17258 15802
rect 1860 15648 1912 15700
rect 5356 15648 5408 15700
rect 5448 15691 5500 15700
rect 5448 15657 5457 15691
rect 5457 15657 5491 15691
rect 5491 15657 5500 15691
rect 5448 15648 5500 15657
rect 5724 15648 5776 15700
rect 2780 15580 2832 15632
rect 3240 15580 3292 15632
rect 3884 15512 3936 15564
rect 4068 15512 4120 15564
rect 204 15444 256 15496
rect 1400 15376 1452 15428
rect 3608 15376 3660 15428
rect 4160 15487 4212 15496
rect 4160 15453 4169 15487
rect 4169 15453 4203 15487
rect 4203 15453 4212 15487
rect 4160 15444 4212 15453
rect 4344 15444 4396 15496
rect 4712 15555 4764 15564
rect 4712 15521 4721 15555
rect 4721 15521 4755 15555
rect 4755 15521 4764 15555
rect 4712 15512 4764 15521
rect 4896 15444 4948 15496
rect 5172 15487 5224 15496
rect 5172 15453 5181 15487
rect 5181 15453 5215 15487
rect 5215 15453 5224 15487
rect 5172 15444 5224 15453
rect 7288 15580 7340 15632
rect 8484 15648 8536 15700
rect 9312 15648 9364 15700
rect 9496 15691 9548 15700
rect 9496 15657 9505 15691
rect 9505 15657 9539 15691
rect 9539 15657 9548 15691
rect 9496 15648 9548 15657
rect 10600 15691 10652 15700
rect 10600 15657 10609 15691
rect 10609 15657 10643 15691
rect 10643 15657 10652 15691
rect 10600 15648 10652 15657
rect 10692 15648 10744 15700
rect 16396 15648 16448 15700
rect 11152 15580 11204 15632
rect 6460 15512 6512 15564
rect 11520 15512 11572 15564
rect 6920 15487 6972 15496
rect 6920 15453 6929 15487
rect 6929 15453 6963 15487
rect 6963 15453 6972 15487
rect 6920 15444 6972 15453
rect 7748 15487 7800 15496
rect 2412 15308 2464 15360
rect 6552 15419 6604 15428
rect 6552 15385 6561 15419
rect 6561 15385 6595 15419
rect 6595 15385 6604 15419
rect 6552 15376 6604 15385
rect 5448 15308 5500 15360
rect 5540 15308 5592 15360
rect 7748 15453 7757 15487
rect 7757 15453 7791 15487
rect 7791 15453 7800 15487
rect 7748 15444 7800 15453
rect 8024 15487 8076 15496
rect 8024 15453 8033 15487
rect 8033 15453 8067 15487
rect 8067 15453 8076 15487
rect 8024 15444 8076 15453
rect 8300 15487 8352 15496
rect 8300 15453 8309 15487
rect 8309 15453 8343 15487
rect 8343 15453 8352 15487
rect 8300 15444 8352 15453
rect 8852 15444 8904 15496
rect 9036 15487 9088 15496
rect 9036 15453 9045 15487
rect 9045 15453 9079 15487
rect 9079 15453 9088 15487
rect 9036 15444 9088 15453
rect 7840 15376 7892 15428
rect 8392 15419 8444 15428
rect 8392 15385 8401 15419
rect 8401 15385 8435 15419
rect 8435 15385 8444 15419
rect 8392 15376 8444 15385
rect 9312 15487 9364 15496
rect 9312 15453 9321 15487
rect 9321 15453 9355 15487
rect 9355 15453 9364 15487
rect 9312 15444 9364 15453
rect 7472 15308 7524 15360
rect 8576 15351 8628 15360
rect 8576 15317 8601 15351
rect 8601 15317 8628 15351
rect 9404 15376 9456 15428
rect 10416 15444 10468 15496
rect 10600 15487 10652 15496
rect 10600 15453 10609 15487
rect 10609 15453 10643 15487
rect 10643 15453 10652 15487
rect 10600 15444 10652 15453
rect 11060 15487 11112 15496
rect 11060 15453 11069 15487
rect 11069 15453 11103 15487
rect 11103 15453 11112 15487
rect 11060 15444 11112 15453
rect 11428 15487 11480 15496
rect 11428 15453 11437 15487
rect 11437 15453 11471 15487
rect 11471 15453 11480 15487
rect 11428 15444 11480 15453
rect 11704 15487 11756 15496
rect 11704 15453 11713 15487
rect 11713 15453 11747 15487
rect 11747 15453 11756 15487
rect 11704 15444 11756 15453
rect 12624 15555 12676 15564
rect 12624 15521 12633 15555
rect 12633 15521 12667 15555
rect 12667 15521 12676 15555
rect 12624 15512 12676 15521
rect 12716 15512 12768 15564
rect 14832 15623 14884 15632
rect 14832 15589 14841 15623
rect 14841 15589 14875 15623
rect 14875 15589 14884 15623
rect 14832 15580 14884 15589
rect 12348 15376 12400 15428
rect 12624 15376 12676 15428
rect 12808 15487 12860 15496
rect 12808 15453 12817 15487
rect 12817 15453 12851 15487
rect 12851 15453 12860 15487
rect 12808 15444 12860 15453
rect 16764 15512 16816 15564
rect 12992 15376 13044 15428
rect 15016 15487 15068 15496
rect 15016 15453 15025 15487
rect 15025 15453 15059 15487
rect 15059 15453 15068 15487
rect 15016 15444 15068 15453
rect 8576 15308 8628 15317
rect 9772 15308 9824 15360
rect 10968 15308 11020 15360
rect 11520 15308 11572 15360
rect 15200 15351 15252 15360
rect 15200 15317 15209 15351
rect 15209 15317 15243 15351
rect 15243 15317 15252 15351
rect 15200 15308 15252 15317
rect 2610 15206 2662 15258
rect 2674 15206 2726 15258
rect 2738 15206 2790 15258
rect 2802 15206 2854 15258
rect 2866 15206 2918 15258
rect 7610 15206 7662 15258
rect 7674 15206 7726 15258
rect 7738 15206 7790 15258
rect 7802 15206 7854 15258
rect 7866 15206 7918 15258
rect 12610 15206 12662 15258
rect 12674 15206 12726 15258
rect 12738 15206 12790 15258
rect 12802 15206 12854 15258
rect 12866 15206 12918 15258
rect 17610 15206 17662 15258
rect 17674 15206 17726 15258
rect 17738 15206 17790 15258
rect 17802 15206 17854 15258
rect 17866 15206 17918 15258
rect 1308 15104 1360 15156
rect 8208 15104 8260 15156
rect 9772 15104 9824 15156
rect 9956 15104 10008 15156
rect 1124 15036 1176 15088
rect 5264 15079 5316 15088
rect 5264 15045 5273 15079
rect 5273 15045 5307 15079
rect 5307 15045 5316 15079
rect 5264 15036 5316 15045
rect 8024 15036 8076 15088
rect 4528 15011 4580 15020
rect 4528 14977 4537 15011
rect 4537 14977 4571 15011
rect 4571 14977 4580 15011
rect 4528 14968 4580 14977
rect 4620 15011 4672 15020
rect 4620 14977 4629 15011
rect 4629 14977 4663 15011
rect 4663 14977 4672 15011
rect 4620 14968 4672 14977
rect 1768 14900 1820 14952
rect 2320 14900 2372 14952
rect 3884 14900 3936 14952
rect 8392 14968 8444 15020
rect 9772 14968 9824 15020
rect 10140 15011 10192 15020
rect 10140 14977 10149 15011
rect 10149 14977 10183 15011
rect 10183 14977 10192 15011
rect 10140 14968 10192 14977
rect 10232 14968 10284 15020
rect 3976 14832 4028 14884
rect 8484 14900 8536 14952
rect 8576 14900 8628 14952
rect 9312 14900 9364 14952
rect 9680 14943 9732 14952
rect 9680 14909 9689 14943
rect 9689 14909 9723 14943
rect 9723 14909 9732 14943
rect 9680 14900 9732 14909
rect 10416 14900 10468 14952
rect 11244 15036 11296 15088
rect 12808 15036 12860 15088
rect 12440 14968 12492 15020
rect 12900 15011 12952 15020
rect 12900 14977 12909 15011
rect 12909 14977 12943 15011
rect 12943 14977 12952 15011
rect 12900 14968 12952 14977
rect 13728 15036 13780 15088
rect 3240 14764 3292 14816
rect 5632 14832 5684 14884
rect 13084 14900 13136 14952
rect 13360 15011 13412 15020
rect 13360 14977 13369 15011
rect 13369 14977 13403 15011
rect 13403 14977 13412 15011
rect 13360 14968 13412 14977
rect 13452 14968 13504 15020
rect 13820 14968 13872 15020
rect 14280 15036 14332 15088
rect 16672 15011 16724 15020
rect 16672 14977 16681 15011
rect 16681 14977 16715 15011
rect 16715 14977 16724 15011
rect 16672 14968 16724 14977
rect 11152 14832 11204 14884
rect 12624 14832 12676 14884
rect 13176 14832 13228 14884
rect 14740 14943 14792 14952
rect 14740 14909 14749 14943
rect 14749 14909 14783 14943
rect 14783 14909 14792 14943
rect 14740 14900 14792 14909
rect 16028 14900 16080 14952
rect 17408 15011 17460 15020
rect 17408 14977 17417 15011
rect 17417 14977 17451 15011
rect 17451 14977 17460 15011
rect 17408 14968 17460 14977
rect 18144 15011 18196 15020
rect 18144 14977 18153 15011
rect 18153 14977 18187 15011
rect 18187 14977 18196 15011
rect 18144 14968 18196 14977
rect 15108 14832 15160 14884
rect 8484 14764 8536 14816
rect 9496 14764 9548 14816
rect 10600 14764 10652 14816
rect 11520 14807 11572 14816
rect 11520 14773 11529 14807
rect 11529 14773 11563 14807
rect 11563 14773 11572 14807
rect 11520 14764 11572 14773
rect 11704 14764 11756 14816
rect 15200 14764 15252 14816
rect 1950 14662 2002 14714
rect 2014 14662 2066 14714
rect 2078 14662 2130 14714
rect 2142 14662 2194 14714
rect 2206 14662 2258 14714
rect 6950 14662 7002 14714
rect 7014 14662 7066 14714
rect 7078 14662 7130 14714
rect 7142 14662 7194 14714
rect 7206 14662 7258 14714
rect 11950 14662 12002 14714
rect 12014 14662 12066 14714
rect 12078 14662 12130 14714
rect 12142 14662 12194 14714
rect 12206 14662 12258 14714
rect 16950 14662 17002 14714
rect 17014 14662 17066 14714
rect 17078 14662 17130 14714
rect 17142 14662 17194 14714
rect 17206 14662 17258 14714
rect 1768 14603 1820 14612
rect 1768 14569 1777 14603
rect 1777 14569 1811 14603
rect 1811 14569 1820 14603
rect 1768 14560 1820 14569
rect 2228 14560 2280 14612
rect 6184 14560 6236 14612
rect 8392 14560 8444 14612
rect 6552 14492 6604 14544
rect 8576 14492 8628 14544
rect 8760 14492 8812 14544
rect 9496 14560 9548 14612
rect 10692 14560 10744 14612
rect 10968 14560 11020 14612
rect 11888 14560 11940 14612
rect 12256 14560 12308 14612
rect 12624 14560 12676 14612
rect 12716 14560 12768 14612
rect 14096 14560 14148 14612
rect 15752 14560 15804 14612
rect 16488 14560 16540 14612
rect 11152 14492 11204 14544
rect 11244 14492 11296 14544
rect 11704 14492 11756 14544
rect 1676 14424 1728 14476
rect 1860 14424 1912 14476
rect 2228 14467 2280 14476
rect 2228 14433 2237 14467
rect 2237 14433 2271 14467
rect 2271 14433 2280 14467
rect 2228 14424 2280 14433
rect 2964 14424 3016 14476
rect 6000 14424 6052 14476
rect 1952 14399 2004 14408
rect 1952 14365 1961 14399
rect 1961 14365 1995 14399
rect 1995 14365 2004 14399
rect 1952 14356 2004 14365
rect 2136 14399 2188 14408
rect 2136 14365 2145 14399
rect 2145 14365 2179 14399
rect 2179 14365 2188 14399
rect 2136 14356 2188 14365
rect 4712 14399 4764 14408
rect 4712 14365 4721 14399
rect 4721 14365 4755 14399
rect 4755 14365 4764 14399
rect 4712 14356 4764 14365
rect 4988 14399 5040 14408
rect 4988 14365 4997 14399
rect 4997 14365 5031 14399
rect 5031 14365 5040 14399
rect 4988 14356 5040 14365
rect 5172 14356 5224 14408
rect 5264 14356 5316 14408
rect 9128 14424 9180 14476
rect 9312 14424 9364 14476
rect 12992 14492 13044 14544
rect 13360 14492 13412 14544
rect 13636 14492 13688 14544
rect 3608 14288 3660 14340
rect 4896 14263 4948 14272
rect 4896 14229 4905 14263
rect 4905 14229 4939 14263
rect 4939 14229 4948 14263
rect 4896 14220 4948 14229
rect 5908 14220 5960 14272
rect 10508 14288 10560 14340
rect 10692 14356 10744 14408
rect 12716 14356 12768 14408
rect 12992 14356 13044 14408
rect 13452 14424 13504 14476
rect 11888 14331 11940 14340
rect 11888 14297 11897 14331
rect 11897 14297 11931 14331
rect 11931 14297 11940 14331
rect 11888 14288 11940 14297
rect 13912 14356 13964 14408
rect 14280 14399 14332 14408
rect 14280 14365 14289 14399
rect 14289 14365 14323 14399
rect 14323 14365 14332 14399
rect 14280 14356 14332 14365
rect 15936 14424 15988 14476
rect 16488 14424 16540 14476
rect 16396 14356 16448 14408
rect 16672 14399 16724 14408
rect 16672 14365 16681 14399
rect 16681 14365 16715 14399
rect 16715 14365 16724 14399
rect 16672 14356 16724 14365
rect 17500 14492 17552 14544
rect 13544 14288 13596 14340
rect 14188 14331 14240 14340
rect 14188 14297 14197 14331
rect 14197 14297 14231 14331
rect 14231 14297 14240 14331
rect 14188 14288 14240 14297
rect 9772 14263 9824 14272
rect 9772 14229 9781 14263
rect 9781 14229 9815 14263
rect 9815 14229 9824 14263
rect 9772 14220 9824 14229
rect 10968 14220 11020 14272
rect 11520 14263 11572 14272
rect 11520 14229 11529 14263
rect 11529 14229 11563 14263
rect 11563 14229 11572 14263
rect 11520 14220 11572 14229
rect 11980 14220 12032 14272
rect 12440 14220 12492 14272
rect 16304 14220 16356 14272
rect 18236 14356 18288 14408
rect 16672 14220 16724 14272
rect 16764 14220 16816 14272
rect 17132 14220 17184 14272
rect 18052 14331 18104 14340
rect 18052 14297 18061 14331
rect 18061 14297 18095 14331
rect 18095 14297 18104 14331
rect 18052 14288 18104 14297
rect 18880 14220 18932 14272
rect 2610 14118 2662 14170
rect 2674 14118 2726 14170
rect 2738 14118 2790 14170
rect 2802 14118 2854 14170
rect 2866 14118 2918 14170
rect 7610 14118 7662 14170
rect 7674 14118 7726 14170
rect 7738 14118 7790 14170
rect 7802 14118 7854 14170
rect 7866 14118 7918 14170
rect 12610 14118 12662 14170
rect 12674 14118 12726 14170
rect 12738 14118 12790 14170
rect 12802 14118 12854 14170
rect 12866 14118 12918 14170
rect 17610 14118 17662 14170
rect 17674 14118 17726 14170
rect 17738 14118 17790 14170
rect 17802 14118 17854 14170
rect 17866 14118 17918 14170
rect 2872 14016 2924 14068
rect 3240 14016 3292 14068
rect 4620 14016 4672 14068
rect 8668 14016 8720 14068
rect 9220 14059 9272 14068
rect 9220 14025 9229 14059
rect 9229 14025 9263 14059
rect 9263 14025 9272 14059
rect 9220 14016 9272 14025
rect 9312 14016 9364 14068
rect 11152 14016 11204 14068
rect 13636 14016 13688 14068
rect 13820 14016 13872 14068
rect 16028 14016 16080 14068
rect 1492 13923 1544 13932
rect 1492 13889 1501 13923
rect 1501 13889 1535 13923
rect 1535 13889 1544 13923
rect 1492 13880 1544 13889
rect 3424 13948 3476 14000
rect 5356 13948 5408 14000
rect 2872 13923 2924 13932
rect 2872 13889 2881 13923
rect 2881 13889 2915 13923
rect 2915 13889 2924 13923
rect 2872 13880 2924 13889
rect 2964 13923 3016 13932
rect 2964 13889 2973 13923
rect 2973 13889 3007 13923
rect 3007 13889 3016 13923
rect 2964 13880 3016 13889
rect 3884 13880 3936 13932
rect 4804 13880 4856 13932
rect 5724 13880 5776 13932
rect 5908 13923 5960 13932
rect 5908 13889 5917 13923
rect 5917 13889 5951 13923
rect 5951 13889 5960 13923
rect 5908 13880 5960 13889
rect 3240 13812 3292 13864
rect 296 13744 348 13796
rect 5172 13812 5224 13864
rect 5356 13812 5408 13864
rect 5540 13812 5592 13864
rect 5816 13812 5868 13864
rect 8116 13948 8168 14000
rect 6368 13923 6420 13932
rect 6368 13889 6377 13923
rect 6377 13889 6411 13923
rect 6411 13889 6420 13923
rect 6368 13880 6420 13889
rect 6460 13923 6512 13932
rect 6460 13889 6469 13923
rect 6469 13889 6503 13923
rect 6503 13889 6512 13923
rect 6460 13880 6512 13889
rect 6644 13923 6696 13932
rect 6644 13889 6653 13923
rect 6653 13889 6687 13923
rect 6687 13889 6696 13923
rect 6644 13880 6696 13889
rect 7748 13880 7800 13932
rect 8024 13880 8076 13932
rect 8668 13880 8720 13932
rect 4988 13744 5040 13796
rect 8484 13812 8536 13864
rect 8944 13923 8996 13932
rect 8944 13889 8953 13923
rect 8953 13889 8987 13923
rect 8987 13889 8996 13923
rect 8944 13880 8996 13889
rect 9312 13880 9364 13932
rect 9128 13812 9180 13864
rect 9220 13847 9272 13864
rect 9220 13813 9229 13847
rect 9229 13813 9263 13847
rect 9263 13813 9272 13847
rect 9220 13812 9272 13813
rect 9588 13812 9640 13864
rect 10968 13812 11020 13864
rect 11612 13812 11664 13864
rect 11704 13812 11756 13864
rect 12440 13880 12492 13932
rect 12716 13880 12768 13932
rect 13912 13948 13964 14000
rect 13176 13880 13228 13932
rect 15752 13880 15804 13932
rect 18236 13923 18288 13932
rect 18236 13889 18245 13923
rect 18245 13889 18279 13923
rect 18279 13889 18288 13923
rect 18236 13880 18288 13889
rect 19340 13880 19392 13932
rect 13728 13812 13780 13864
rect 16580 13812 16632 13864
rect 6736 13744 6788 13796
rect 3608 13676 3660 13728
rect 3976 13676 4028 13728
rect 5172 13676 5224 13728
rect 5724 13719 5776 13728
rect 5724 13685 5733 13719
rect 5733 13685 5767 13719
rect 5767 13685 5776 13719
rect 5724 13676 5776 13685
rect 6276 13676 6328 13728
rect 6828 13676 6880 13728
rect 7564 13676 7616 13728
rect 7932 13676 7984 13728
rect 8484 13676 8536 13728
rect 14556 13744 14608 13796
rect 10416 13676 10468 13728
rect 11428 13676 11480 13728
rect 12256 13676 12308 13728
rect 12440 13676 12492 13728
rect 12532 13676 12584 13728
rect 12716 13676 12768 13728
rect 13452 13676 13504 13728
rect 14924 13676 14976 13728
rect 17132 13676 17184 13728
rect 1950 13574 2002 13626
rect 2014 13574 2066 13626
rect 2078 13574 2130 13626
rect 2142 13574 2194 13626
rect 2206 13574 2258 13626
rect 6950 13574 7002 13626
rect 7014 13574 7066 13626
rect 7078 13574 7130 13626
rect 7142 13574 7194 13626
rect 7206 13574 7258 13626
rect 11950 13574 12002 13626
rect 12014 13574 12066 13626
rect 12078 13574 12130 13626
rect 12142 13574 12194 13626
rect 12206 13574 12258 13626
rect 16950 13574 17002 13626
rect 17014 13574 17066 13626
rect 17078 13574 17130 13626
rect 17142 13574 17194 13626
rect 17206 13574 17258 13626
rect 2228 13472 2280 13524
rect 3148 13515 3200 13524
rect 3148 13481 3157 13515
rect 3157 13481 3191 13515
rect 3191 13481 3200 13515
rect 3148 13472 3200 13481
rect 4712 13472 4764 13524
rect 4988 13472 5040 13524
rect 5356 13472 5408 13524
rect 5448 13472 5500 13524
rect 9036 13472 9088 13524
rect 9496 13515 9548 13524
rect 9496 13481 9505 13515
rect 9505 13481 9539 13515
rect 9539 13481 9548 13515
rect 9496 13472 9548 13481
rect 10048 13472 10100 13524
rect 17224 13472 17276 13524
rect 18420 13515 18472 13524
rect 18420 13481 18429 13515
rect 18429 13481 18463 13515
rect 18463 13481 18472 13515
rect 18420 13472 18472 13481
rect 6736 13404 6788 13456
rect 940 13336 992 13388
rect 5172 13336 5224 13388
rect 5448 13336 5500 13388
rect 6092 13336 6144 13388
rect 6460 13336 6512 13388
rect 6920 13336 6972 13388
rect 2320 13268 2372 13320
rect 2504 13311 2556 13320
rect 2504 13277 2513 13311
rect 2513 13277 2547 13311
rect 2547 13277 2556 13311
rect 2504 13268 2556 13277
rect 2596 13311 2648 13320
rect 2596 13277 2605 13311
rect 2605 13277 2639 13311
rect 2639 13277 2648 13311
rect 2596 13268 2648 13277
rect 2872 13311 2924 13320
rect 2872 13277 2881 13311
rect 2881 13277 2915 13311
rect 2915 13277 2924 13311
rect 2872 13268 2924 13277
rect 2964 13311 3016 13320
rect 2964 13277 2973 13311
rect 2973 13277 3007 13311
rect 3007 13277 3016 13311
rect 2964 13268 3016 13277
rect 3148 13268 3200 13320
rect 4068 13268 4120 13320
rect 4528 13268 4580 13320
rect 6276 13311 6328 13320
rect 6276 13277 6285 13311
rect 6285 13277 6319 13311
rect 6319 13277 6328 13311
rect 6276 13268 6328 13277
rect 8208 13404 8260 13456
rect 10232 13404 10284 13456
rect 11060 13404 11112 13456
rect 7288 13336 7340 13388
rect 8116 13336 8168 13388
rect 9312 13336 9364 13388
rect 1768 13132 1820 13184
rect 3792 13200 3844 13252
rect 4252 13200 4304 13252
rect 5356 13200 5408 13252
rect 6092 13200 6144 13252
rect 7932 13268 7984 13320
rect 8300 13268 8352 13320
rect 9864 13336 9916 13388
rect 10876 13336 10928 13388
rect 11888 13336 11940 13388
rect 11980 13336 12032 13388
rect 12440 13336 12492 13388
rect 19432 13404 19484 13456
rect 14004 13336 14056 13388
rect 11244 13311 11296 13320
rect 11244 13277 11253 13311
rect 11253 13277 11287 13311
rect 11287 13277 11296 13311
rect 11244 13268 11296 13277
rect 12624 13311 12676 13320
rect 12624 13277 12633 13311
rect 12633 13277 12667 13311
rect 12667 13277 12676 13311
rect 12624 13268 12676 13277
rect 8208 13200 8260 13252
rect 9864 13200 9916 13252
rect 7012 13132 7064 13184
rect 11796 13200 11848 13252
rect 13084 13268 13136 13320
rect 13268 13268 13320 13320
rect 13636 13268 13688 13320
rect 14648 13268 14700 13320
rect 15200 13268 15252 13320
rect 15476 13311 15528 13320
rect 15476 13277 15485 13311
rect 15485 13277 15519 13311
rect 15519 13277 15528 13311
rect 15476 13268 15528 13277
rect 16672 13268 16724 13320
rect 16856 13200 16908 13252
rect 17500 13200 17552 13252
rect 18236 13311 18288 13320
rect 18236 13277 18245 13311
rect 18245 13277 18279 13311
rect 18279 13277 18288 13311
rect 18236 13268 18288 13277
rect 11612 13175 11664 13184
rect 11612 13141 11621 13175
rect 11621 13141 11655 13175
rect 11655 13141 11664 13175
rect 11612 13132 11664 13141
rect 11704 13132 11756 13184
rect 15844 13132 15896 13184
rect 2610 13030 2662 13082
rect 2674 13030 2726 13082
rect 2738 13030 2790 13082
rect 2802 13030 2854 13082
rect 2866 13030 2918 13082
rect 7610 13030 7662 13082
rect 7674 13030 7726 13082
rect 7738 13030 7790 13082
rect 7802 13030 7854 13082
rect 7866 13030 7918 13082
rect 12610 13030 12662 13082
rect 12674 13030 12726 13082
rect 12738 13030 12790 13082
rect 12802 13030 12854 13082
rect 12866 13030 12918 13082
rect 17610 13030 17662 13082
rect 17674 13030 17726 13082
rect 17738 13030 17790 13082
rect 17802 13030 17854 13082
rect 17866 13030 17918 13082
rect 2320 12928 2372 12980
rect 2688 12928 2740 12980
rect 2964 12928 3016 12980
rect 7380 12928 7432 12980
rect 7656 12928 7708 12980
rect 9220 12928 9272 12980
rect 11520 12928 11572 12980
rect 11888 12928 11940 12980
rect 15016 12928 15068 12980
rect 15292 12928 15344 12980
rect 15476 12928 15528 12980
rect 16028 12928 16080 12980
rect 18052 12928 18104 12980
rect 1952 12860 2004 12912
rect 2228 12860 2280 12912
rect 3516 12860 3568 12912
rect 4712 12860 4764 12912
rect 4988 12903 5040 12912
rect 4988 12869 4997 12903
rect 4997 12869 5031 12903
rect 5031 12869 5040 12903
rect 4988 12860 5040 12869
rect 2780 12792 2832 12844
rect 3056 12835 3108 12844
rect 3056 12801 3065 12835
rect 3065 12801 3099 12835
rect 3099 12801 3108 12835
rect 3056 12792 3108 12801
rect 3240 12835 3292 12844
rect 3240 12801 3249 12835
rect 3249 12801 3283 12835
rect 3283 12801 3292 12835
rect 3240 12792 3292 12801
rect 480 12724 532 12776
rect 1860 12724 1912 12776
rect 2504 12767 2556 12776
rect 2504 12733 2513 12767
rect 2513 12733 2547 12767
rect 2547 12733 2556 12767
rect 2504 12724 2556 12733
rect 2964 12767 3016 12776
rect 2964 12733 2973 12767
rect 2973 12733 3007 12767
rect 3007 12733 3016 12767
rect 2964 12724 3016 12733
rect 4620 12835 4672 12844
rect 4620 12801 4629 12835
rect 4629 12801 4663 12835
rect 4663 12801 4672 12835
rect 4620 12792 4672 12801
rect 10416 12860 10468 12912
rect 5356 12835 5408 12844
rect 5356 12801 5365 12835
rect 5365 12801 5399 12835
rect 5399 12801 5408 12835
rect 5356 12792 5408 12801
rect 5448 12835 5500 12844
rect 5448 12801 5457 12835
rect 5457 12801 5491 12835
rect 5491 12801 5500 12835
rect 5448 12792 5500 12801
rect 5632 12792 5684 12844
rect 6552 12792 6604 12844
rect 6736 12835 6788 12844
rect 6736 12801 6745 12835
rect 6745 12801 6779 12835
rect 6779 12801 6788 12835
rect 6736 12792 6788 12801
rect 7012 12835 7064 12844
rect 7012 12801 7021 12835
rect 7021 12801 7055 12835
rect 7055 12801 7064 12835
rect 7012 12792 7064 12801
rect 7564 12835 7616 12844
rect 7564 12801 7576 12835
rect 7576 12801 7610 12835
rect 7610 12801 7616 12835
rect 7564 12792 7616 12801
rect 7748 12792 7800 12844
rect 8392 12792 8444 12844
rect 9312 12792 9364 12844
rect 8300 12724 8352 12776
rect 9036 12724 9088 12776
rect 9772 12724 9824 12776
rect 10048 12835 10100 12844
rect 10048 12801 10057 12835
rect 10057 12801 10091 12835
rect 10091 12801 10100 12835
rect 10048 12792 10100 12801
rect 13084 12860 13136 12912
rect 13268 12860 13320 12912
rect 10876 12792 10928 12844
rect 10968 12835 11020 12844
rect 10968 12801 10977 12835
rect 10977 12801 11011 12835
rect 11011 12801 11020 12835
rect 10968 12792 11020 12801
rect 11244 12792 11296 12844
rect 11336 12792 11388 12844
rect 11980 12835 12032 12844
rect 11980 12801 11989 12835
rect 11989 12801 12023 12835
rect 12023 12801 12032 12835
rect 11980 12792 12032 12801
rect 12072 12792 12124 12844
rect 10416 12724 10468 12776
rect 3240 12588 3292 12640
rect 3608 12631 3660 12640
rect 3608 12597 3617 12631
rect 3617 12597 3651 12631
rect 3651 12597 3660 12631
rect 3608 12588 3660 12597
rect 3884 12631 3936 12640
rect 3884 12597 3893 12631
rect 3893 12597 3927 12631
rect 3927 12597 3936 12631
rect 3884 12588 3936 12597
rect 4620 12656 4672 12708
rect 7564 12656 7616 12708
rect 7748 12656 7800 12708
rect 9588 12656 9640 12708
rect 9956 12656 10008 12708
rect 11704 12724 11756 12776
rect 11796 12724 11848 12776
rect 12256 12724 12308 12776
rect 12440 12792 12492 12844
rect 12900 12792 12952 12844
rect 13452 12792 13504 12844
rect 14832 12792 14884 12844
rect 15016 12792 15068 12844
rect 16028 12835 16080 12844
rect 12716 12724 12768 12776
rect 13912 12724 13964 12776
rect 16028 12801 16037 12835
rect 16037 12801 16071 12835
rect 16071 12801 16080 12835
rect 16028 12792 16080 12801
rect 16304 12860 16356 12912
rect 15936 12724 15988 12776
rect 10600 12699 10652 12708
rect 10600 12665 10609 12699
rect 10609 12665 10643 12699
rect 10643 12665 10652 12699
rect 10600 12656 10652 12665
rect 6736 12588 6788 12640
rect 6828 12588 6880 12640
rect 7012 12588 7064 12640
rect 8392 12588 8444 12640
rect 10508 12588 10560 12640
rect 10692 12588 10744 12640
rect 11152 12588 11204 12640
rect 11244 12588 11296 12640
rect 13176 12656 13228 12708
rect 13452 12656 13504 12708
rect 17224 12792 17276 12844
rect 17684 12835 17736 12844
rect 17684 12801 17693 12835
rect 17693 12801 17727 12835
rect 17727 12801 17736 12835
rect 17684 12792 17736 12801
rect 18328 12860 18380 12912
rect 18236 12724 18288 12776
rect 12624 12588 12676 12640
rect 13544 12588 13596 12640
rect 14188 12588 14240 12640
rect 17408 12588 17460 12640
rect 18512 12588 18564 12640
rect 1950 12486 2002 12538
rect 2014 12486 2066 12538
rect 2078 12486 2130 12538
rect 2142 12486 2194 12538
rect 2206 12486 2258 12538
rect 6950 12486 7002 12538
rect 7014 12486 7066 12538
rect 7078 12486 7130 12538
rect 7142 12486 7194 12538
rect 7206 12486 7258 12538
rect 11950 12486 12002 12538
rect 12014 12486 12066 12538
rect 12078 12486 12130 12538
rect 12142 12486 12194 12538
rect 12206 12486 12258 12538
rect 16950 12486 17002 12538
rect 17014 12486 17066 12538
rect 17078 12486 17130 12538
rect 17142 12486 17194 12538
rect 17206 12486 17258 12538
rect 2136 12384 2188 12436
rect 3792 12384 3844 12436
rect 4160 12384 4212 12436
rect 5632 12384 5684 12436
rect 5816 12384 5868 12436
rect 7656 12384 7708 12436
rect 8208 12384 8260 12436
rect 9036 12384 9088 12436
rect 9772 12384 9824 12436
rect 10140 12384 10192 12436
rect 12992 12384 13044 12436
rect 13544 12384 13596 12436
rect 14832 12384 14884 12436
rect 15108 12384 15160 12436
rect 16212 12384 16264 12436
rect 8116 12316 8168 12368
rect 8944 12316 8996 12368
rect 9680 12316 9732 12368
rect 10324 12316 10376 12368
rect 11244 12316 11296 12368
rect 11336 12316 11388 12368
rect 14648 12316 14700 12368
rect 15752 12316 15804 12368
rect 16488 12316 16540 12368
rect 17500 12384 17552 12436
rect 18144 12316 18196 12368
rect 1308 12248 1360 12300
rect 3700 12248 3752 12300
rect 5908 12291 5960 12300
rect 5908 12257 5917 12291
rect 5917 12257 5951 12291
rect 5951 12257 5960 12291
rect 5908 12248 5960 12257
rect 6000 12248 6052 12300
rect 7012 12248 7064 12300
rect 7288 12248 7340 12300
rect 1400 12180 1452 12232
rect 2688 12112 2740 12164
rect 3332 12112 3384 12164
rect 3700 12112 3752 12164
rect 4252 12223 4304 12232
rect 4252 12189 4261 12223
rect 4261 12189 4295 12223
rect 4295 12189 4304 12223
rect 4252 12180 4304 12189
rect 4436 12180 4488 12232
rect 4988 12180 5040 12232
rect 5448 12180 5500 12232
rect 6184 12180 6236 12232
rect 5632 12112 5684 12164
rect 6552 12112 6604 12164
rect 7380 12112 7432 12164
rect 8760 12112 8812 12164
rect 9220 12223 9272 12232
rect 9220 12189 9229 12223
rect 9229 12189 9263 12223
rect 9263 12189 9272 12223
rect 9220 12180 9272 12189
rect 9312 12112 9364 12164
rect 3516 12044 3568 12096
rect 10232 12180 10284 12232
rect 10692 12180 10744 12232
rect 11612 12248 11664 12300
rect 12440 12248 12492 12300
rect 12624 12180 12676 12232
rect 13084 12248 13136 12300
rect 13544 12248 13596 12300
rect 12992 12223 13044 12232
rect 12992 12189 13001 12223
rect 13001 12189 13035 12223
rect 13035 12189 13044 12223
rect 12992 12180 13044 12189
rect 13176 12223 13228 12232
rect 13176 12189 13185 12223
rect 13185 12189 13219 12223
rect 13219 12189 13228 12223
rect 13176 12180 13228 12189
rect 9588 12112 9640 12164
rect 16948 12248 17000 12300
rect 17408 12291 17460 12300
rect 17408 12257 17417 12291
rect 17417 12257 17451 12291
rect 17451 12257 17460 12291
rect 17408 12248 17460 12257
rect 14004 12112 14056 12164
rect 9772 12044 9824 12096
rect 10784 12044 10836 12096
rect 12256 12044 12308 12096
rect 12716 12044 12768 12096
rect 13176 12044 13228 12096
rect 13360 12044 13412 12096
rect 14280 12112 14332 12164
rect 15384 12180 15436 12232
rect 16304 12223 16356 12232
rect 16304 12189 16313 12223
rect 16313 12189 16347 12223
rect 16347 12189 16356 12223
rect 16304 12180 16356 12189
rect 16488 12223 16540 12232
rect 16488 12189 16497 12223
rect 16497 12189 16531 12223
rect 16531 12189 16540 12223
rect 16488 12180 16540 12189
rect 15292 12112 15344 12164
rect 15936 12112 15988 12164
rect 16672 12180 16724 12232
rect 17040 12223 17092 12232
rect 17040 12189 17049 12223
rect 17049 12189 17083 12223
rect 17083 12189 17092 12223
rect 17040 12180 17092 12189
rect 14556 12044 14608 12096
rect 14648 12044 14700 12096
rect 18144 12223 18196 12232
rect 18144 12189 18153 12223
rect 18153 12189 18187 12223
rect 18187 12189 18196 12223
rect 18144 12180 18196 12189
rect 18972 12180 19024 12232
rect 18604 12112 18656 12164
rect 18144 12044 18196 12096
rect 19248 12044 19300 12096
rect 2610 11942 2662 11994
rect 2674 11942 2726 11994
rect 2738 11942 2790 11994
rect 2802 11942 2854 11994
rect 2866 11942 2918 11994
rect 7610 11942 7662 11994
rect 7674 11942 7726 11994
rect 7738 11942 7790 11994
rect 7802 11942 7854 11994
rect 7866 11942 7918 11994
rect 12610 11942 12662 11994
rect 12674 11942 12726 11994
rect 12738 11942 12790 11994
rect 12802 11942 12854 11994
rect 12866 11942 12918 11994
rect 17610 11942 17662 11994
rect 17674 11942 17726 11994
rect 17738 11942 17790 11994
rect 17802 11942 17854 11994
rect 17866 11942 17918 11994
rect 2504 11840 2556 11892
rect 4068 11840 4120 11892
rect 5264 11840 5316 11892
rect 5448 11840 5500 11892
rect 3424 11772 3476 11824
rect 3884 11772 3936 11824
rect 6368 11772 6420 11824
rect 7380 11883 7432 11892
rect 7380 11849 7389 11883
rect 7389 11849 7423 11883
rect 7423 11849 7432 11883
rect 7380 11840 7432 11849
rect 7564 11840 7616 11892
rect 9772 11840 9824 11892
rect 3056 11747 3108 11756
rect 3056 11713 3065 11747
rect 3065 11713 3099 11747
rect 3099 11713 3108 11747
rect 3056 11704 3108 11713
rect 3608 11704 3660 11756
rect 4160 11704 4212 11756
rect 4436 11704 4488 11756
rect 5172 11747 5224 11756
rect 5172 11713 5181 11747
rect 5181 11713 5215 11747
rect 5215 11713 5224 11747
rect 5172 11704 5224 11713
rect 7288 11772 7340 11824
rect 10140 11840 10192 11892
rect 3516 11679 3568 11688
rect 3516 11645 3525 11679
rect 3525 11645 3559 11679
rect 3559 11645 3568 11679
rect 3516 11636 3568 11645
rect 4252 11636 4304 11688
rect 2596 11568 2648 11620
rect 572 11500 624 11552
rect 1492 11500 1544 11552
rect 1860 11500 1912 11552
rect 2136 11500 2188 11552
rect 2504 11500 2556 11552
rect 2872 11500 2924 11552
rect 4712 11500 4764 11552
rect 7012 11747 7064 11756
rect 7012 11713 7021 11747
rect 7021 11713 7055 11747
rect 7055 11713 7064 11747
rect 7012 11704 7064 11713
rect 7380 11704 7432 11756
rect 10048 11772 10100 11824
rect 12808 11840 12860 11892
rect 13360 11840 13412 11892
rect 13912 11840 13964 11892
rect 16488 11840 16540 11892
rect 17040 11840 17092 11892
rect 10876 11772 10928 11824
rect 11060 11772 11112 11824
rect 13728 11772 13780 11824
rect 15476 11772 15528 11824
rect 16580 11772 16632 11824
rect 16856 11772 16908 11824
rect 6092 11568 6144 11620
rect 6460 11568 6512 11620
rect 6552 11568 6604 11620
rect 6736 11568 6788 11620
rect 7748 11747 7800 11756
rect 7748 11713 7757 11747
rect 7757 11713 7791 11747
rect 7791 11713 7800 11747
rect 7748 11704 7800 11713
rect 8392 11704 8444 11756
rect 9496 11704 9548 11756
rect 9680 11704 9732 11756
rect 7840 11636 7892 11688
rect 8024 11679 8076 11688
rect 8024 11645 8033 11679
rect 8033 11645 8067 11679
rect 8067 11645 8076 11679
rect 8024 11636 8076 11645
rect 5540 11500 5592 11552
rect 5724 11500 5776 11552
rect 6368 11543 6420 11552
rect 6368 11509 6377 11543
rect 6377 11509 6411 11543
rect 6411 11509 6420 11543
rect 6368 11500 6420 11509
rect 8392 11568 8444 11620
rect 9956 11636 10008 11688
rect 10508 11704 10560 11756
rect 10784 11704 10836 11756
rect 11152 11747 11204 11756
rect 11152 11713 11161 11747
rect 11161 11713 11195 11747
rect 11195 11713 11204 11747
rect 11152 11704 11204 11713
rect 11520 11704 11572 11756
rect 12808 11704 12860 11756
rect 17408 11747 17460 11756
rect 17408 11713 17417 11747
rect 17417 11713 17451 11747
rect 17451 11713 17460 11747
rect 17408 11704 17460 11713
rect 18236 11815 18288 11824
rect 18236 11781 18245 11815
rect 18245 11781 18279 11815
rect 18279 11781 18288 11815
rect 18236 11772 18288 11781
rect 8944 11568 8996 11620
rect 10048 11568 10100 11620
rect 11428 11568 11480 11620
rect 11796 11568 11848 11620
rect 12348 11636 12400 11688
rect 14004 11636 14056 11688
rect 14372 11679 14424 11688
rect 14372 11645 14381 11679
rect 14381 11645 14415 11679
rect 14415 11645 14424 11679
rect 14372 11636 14424 11645
rect 13268 11568 13320 11620
rect 14648 11679 14700 11688
rect 14648 11645 14657 11679
rect 14657 11645 14691 11679
rect 14691 11645 14700 11679
rect 14648 11636 14700 11645
rect 15936 11636 15988 11688
rect 16764 11636 16816 11688
rect 18512 11636 18564 11688
rect 14832 11568 14884 11620
rect 7932 11500 7984 11552
rect 8576 11500 8628 11552
rect 13728 11500 13780 11552
rect 15844 11500 15896 11552
rect 16764 11500 16816 11552
rect 17500 11500 17552 11552
rect 1950 11398 2002 11450
rect 2014 11398 2066 11450
rect 2078 11398 2130 11450
rect 2142 11398 2194 11450
rect 2206 11398 2258 11450
rect 6950 11398 7002 11450
rect 7014 11398 7066 11450
rect 7078 11398 7130 11450
rect 7142 11398 7194 11450
rect 7206 11398 7258 11450
rect 11950 11398 12002 11450
rect 12014 11398 12066 11450
rect 12078 11398 12130 11450
rect 12142 11398 12194 11450
rect 12206 11398 12258 11450
rect 16950 11398 17002 11450
rect 17014 11398 17066 11450
rect 17078 11398 17130 11450
rect 17142 11398 17194 11450
rect 17206 11398 17258 11450
rect 1400 11296 1452 11348
rect 2228 11296 2280 11348
rect 2596 11296 2648 11348
rect 3700 11296 3752 11348
rect 4160 11296 4212 11348
rect 4620 11296 4672 11348
rect 1584 11228 1636 11280
rect 2964 11228 3016 11280
rect 4068 11228 4120 11280
rect 4436 11228 4488 11280
rect 1492 11160 1544 11212
rect 1768 11160 1820 11212
rect 4620 11160 4672 11212
rect 6000 11296 6052 11348
rect 6736 11296 6788 11348
rect 7104 11296 7156 11348
rect 1400 11135 1452 11144
rect 1400 11101 1409 11135
rect 1409 11101 1443 11135
rect 1443 11101 1452 11135
rect 1400 11092 1452 11101
rect 3884 11092 3936 11144
rect 8116 11228 8168 11280
rect 10876 11296 10928 11348
rect 14188 11296 14240 11348
rect 14740 11296 14792 11348
rect 16948 11296 17000 11348
rect 10784 11228 10836 11280
rect 5724 11160 5776 11212
rect 5080 11135 5132 11144
rect 5080 11101 5089 11135
rect 5089 11101 5123 11135
rect 5123 11101 5132 11135
rect 5080 11092 5132 11101
rect 1768 11024 1820 11076
rect 3056 11024 3108 11076
rect 4804 11024 4856 11076
rect 5448 11092 5500 11144
rect 6000 11135 6052 11144
rect 6000 11101 6009 11135
rect 6009 11101 6043 11135
rect 6043 11101 6052 11135
rect 6000 11092 6052 11101
rect 6184 11135 6236 11144
rect 6184 11101 6201 11135
rect 6201 11101 6235 11135
rect 6235 11101 6236 11135
rect 6920 11160 6972 11212
rect 7104 11160 7156 11212
rect 7472 11160 7524 11212
rect 8576 11160 8628 11212
rect 8760 11160 8812 11212
rect 9496 11160 9548 11212
rect 10324 11160 10376 11212
rect 6184 11092 6236 11101
rect 6828 11092 6880 11144
rect 1400 10956 1452 11008
rect 3424 10956 3476 11008
rect 6736 10956 6788 11008
rect 7012 11024 7064 11076
rect 7748 11024 7800 11076
rect 7840 11024 7892 11076
rect 8944 11024 8996 11076
rect 9220 11067 9272 11076
rect 9220 11033 9229 11067
rect 9229 11033 9263 11067
rect 9263 11033 9272 11067
rect 9220 11024 9272 11033
rect 10048 11135 10100 11144
rect 10048 11101 10057 11135
rect 10057 11101 10091 11135
rect 10091 11101 10100 11135
rect 10048 11092 10100 11101
rect 10968 11135 11020 11144
rect 10968 11101 10977 11135
rect 10977 11101 11011 11135
rect 11011 11101 11020 11135
rect 10968 11092 11020 11101
rect 11244 11160 11296 11212
rect 12532 11160 12584 11212
rect 12716 11228 12768 11280
rect 13820 11228 13872 11280
rect 15844 11271 15896 11280
rect 15844 11237 15853 11271
rect 15853 11237 15887 11271
rect 15887 11237 15896 11271
rect 15844 11228 15896 11237
rect 17960 11228 18012 11280
rect 11704 11092 11756 11144
rect 11888 11092 11940 11144
rect 12716 11092 12768 11144
rect 13176 11092 13228 11144
rect 14372 11092 14424 11144
rect 15660 11092 15712 11144
rect 15844 11092 15896 11144
rect 16856 11203 16908 11212
rect 16856 11169 16865 11203
rect 16865 11169 16899 11203
rect 16899 11169 16908 11203
rect 16856 11160 16908 11169
rect 9496 10956 9548 11008
rect 10048 10956 10100 11008
rect 11612 10956 11664 11008
rect 11980 11024 12032 11076
rect 12440 11024 12492 11076
rect 16488 11024 16540 11076
rect 17500 11135 17552 11144
rect 17500 11101 17509 11135
rect 17509 11101 17543 11135
rect 17543 11101 17552 11135
rect 17500 11092 17552 11101
rect 17776 11135 17828 11144
rect 17776 11101 17785 11135
rect 17785 11101 17819 11135
rect 17819 11101 17828 11135
rect 17776 11092 17828 11101
rect 18052 11092 18104 11144
rect 17408 11024 17460 11076
rect 12164 10956 12216 11008
rect 15108 10956 15160 11008
rect 15568 10956 15620 11008
rect 17868 10956 17920 11008
rect 18696 10956 18748 11008
rect 2610 10854 2662 10906
rect 2674 10854 2726 10906
rect 2738 10854 2790 10906
rect 2802 10854 2854 10906
rect 2866 10854 2918 10906
rect 7610 10854 7662 10906
rect 7674 10854 7726 10906
rect 7738 10854 7790 10906
rect 7802 10854 7854 10906
rect 7866 10854 7918 10906
rect 12610 10854 12662 10906
rect 12674 10854 12726 10906
rect 12738 10854 12790 10906
rect 12802 10854 12854 10906
rect 12866 10854 12918 10906
rect 17610 10854 17662 10906
rect 17674 10854 17726 10906
rect 17738 10854 17790 10906
rect 17802 10854 17854 10906
rect 17866 10854 17918 10906
rect 2228 10752 2280 10804
rect 2596 10752 2648 10804
rect 3424 10752 3476 10804
rect 3608 10752 3660 10804
rect 4344 10752 4396 10804
rect 4896 10752 4948 10804
rect 4988 10752 5040 10804
rect 5356 10752 5408 10804
rect 5448 10752 5500 10804
rect 8208 10752 8260 10804
rect 2872 10684 2924 10736
rect 4712 10684 4764 10736
rect 4804 10684 4856 10736
rect 3608 10616 3660 10668
rect 3976 10659 4028 10668
rect 3976 10625 3985 10659
rect 3985 10625 4019 10659
rect 4019 10625 4028 10659
rect 3976 10616 4028 10625
rect 4344 10616 4396 10668
rect 4252 10548 4304 10600
rect 5172 10548 5224 10600
rect 5264 10548 5316 10600
rect 5448 10591 5500 10600
rect 5448 10557 5457 10591
rect 5457 10557 5491 10591
rect 5491 10557 5500 10591
rect 5448 10548 5500 10557
rect 6000 10616 6052 10668
rect 6092 10548 6144 10600
rect 6276 10616 6328 10668
rect 6828 10616 6880 10668
rect 7840 10684 7892 10736
rect 11796 10752 11848 10804
rect 12624 10752 12676 10804
rect 13268 10752 13320 10804
rect 13636 10752 13688 10804
rect 14188 10752 14240 10804
rect 7196 10659 7248 10668
rect 7196 10625 7205 10659
rect 7205 10625 7239 10659
rect 7239 10625 7248 10659
rect 7196 10616 7248 10625
rect 7288 10659 7340 10668
rect 7288 10625 7297 10659
rect 7297 10625 7331 10659
rect 7331 10625 7340 10659
rect 7288 10616 7340 10625
rect 7656 10616 7708 10668
rect 9496 10684 9548 10736
rect 9772 10684 9824 10736
rect 9956 10684 10008 10736
rect 11888 10684 11940 10736
rect 8208 10616 8260 10668
rect 11060 10616 11112 10668
rect 7472 10548 7524 10600
rect 7748 10548 7800 10600
rect 11520 10616 11572 10668
rect 11612 10659 11664 10668
rect 11612 10625 11621 10659
rect 11621 10625 11655 10659
rect 11655 10625 11664 10659
rect 11612 10616 11664 10625
rect 11796 10659 11848 10668
rect 11796 10625 11805 10659
rect 11805 10625 11839 10659
rect 11839 10625 11848 10659
rect 11796 10616 11848 10625
rect 12164 10616 12216 10668
rect 12716 10616 12768 10668
rect 12900 10616 12952 10668
rect 3976 10480 4028 10532
rect 5908 10480 5960 10532
rect 6000 10523 6052 10532
rect 6000 10489 6009 10523
rect 6009 10489 6043 10523
rect 6043 10489 6052 10523
rect 6000 10480 6052 10489
rect 3516 10412 3568 10464
rect 3700 10412 3752 10464
rect 5724 10412 5776 10464
rect 7104 10480 7156 10532
rect 12072 10548 12124 10600
rect 12808 10548 12860 10600
rect 13544 10548 13596 10600
rect 14004 10659 14056 10668
rect 14004 10625 14013 10659
rect 14013 10625 14047 10659
rect 14047 10625 14056 10659
rect 14004 10616 14056 10625
rect 14188 10616 14240 10668
rect 15108 10752 15160 10804
rect 15476 10752 15528 10804
rect 14832 10684 14884 10736
rect 15660 10752 15712 10804
rect 17776 10752 17828 10804
rect 18420 10752 18472 10804
rect 15108 10659 15160 10668
rect 15108 10625 15117 10659
rect 15117 10625 15151 10659
rect 15151 10625 15160 10659
rect 15108 10616 15160 10625
rect 15568 10616 15620 10668
rect 16212 10616 16264 10668
rect 16948 10684 17000 10736
rect 14464 10548 14516 10600
rect 14832 10548 14884 10600
rect 11520 10480 11572 10532
rect 11796 10480 11848 10532
rect 14004 10480 14056 10532
rect 14556 10480 14608 10532
rect 17500 10616 17552 10668
rect 17960 10727 18012 10736
rect 17960 10693 17969 10727
rect 17969 10693 18003 10727
rect 18003 10693 18012 10727
rect 17960 10684 18012 10693
rect 18052 10616 18104 10668
rect 19156 10616 19208 10668
rect 17040 10548 17092 10600
rect 6460 10455 6512 10464
rect 6460 10421 6469 10455
rect 6469 10421 6503 10455
rect 6503 10421 6512 10455
rect 6460 10412 6512 10421
rect 6552 10412 6604 10464
rect 7656 10412 7708 10464
rect 8024 10412 8076 10464
rect 8300 10412 8352 10464
rect 10784 10412 10836 10464
rect 10968 10412 11020 10464
rect 13268 10412 13320 10464
rect 13912 10412 13964 10464
rect 17500 10523 17552 10532
rect 17500 10489 17509 10523
rect 17509 10489 17543 10523
rect 17543 10489 17552 10523
rect 17500 10480 17552 10489
rect 15384 10455 15436 10464
rect 15384 10421 15393 10455
rect 15393 10421 15427 10455
rect 15427 10421 15436 10455
rect 15384 10412 15436 10421
rect 15844 10412 15896 10464
rect 16304 10412 16356 10464
rect 17040 10412 17092 10464
rect 17868 10412 17920 10464
rect 18144 10412 18196 10464
rect 1950 10310 2002 10362
rect 2014 10310 2066 10362
rect 2078 10310 2130 10362
rect 2142 10310 2194 10362
rect 2206 10310 2258 10362
rect 6950 10310 7002 10362
rect 7014 10310 7066 10362
rect 7078 10310 7130 10362
rect 7142 10310 7194 10362
rect 7206 10310 7258 10362
rect 11950 10310 12002 10362
rect 12014 10310 12066 10362
rect 12078 10310 12130 10362
rect 12142 10310 12194 10362
rect 12206 10310 12258 10362
rect 16950 10310 17002 10362
rect 17014 10310 17066 10362
rect 17078 10310 17130 10362
rect 17142 10310 17194 10362
rect 17206 10310 17258 10362
rect 1400 10208 1452 10260
rect 1952 10208 2004 10260
rect 3976 10208 4028 10260
rect 4344 10208 4396 10260
rect 4988 10208 5040 10260
rect 1860 10140 1912 10192
rect 2136 10140 2188 10192
rect 2228 10140 2280 10192
rect 2596 10140 2648 10192
rect 1676 10072 1728 10124
rect 1216 10004 1268 10056
rect 1400 10004 1452 10056
rect 2872 10072 2924 10124
rect 3056 10047 3108 10056
rect 3056 10013 3065 10047
rect 3065 10013 3099 10047
rect 3099 10013 3108 10047
rect 3056 10004 3108 10013
rect 3884 10140 3936 10192
rect 5356 10140 5408 10192
rect 6368 10072 6420 10124
rect 2688 9936 2740 9988
rect 3608 10004 3660 10056
rect 4252 10047 4304 10056
rect 4252 10013 4261 10047
rect 4261 10013 4295 10047
rect 4295 10013 4304 10047
rect 4252 10004 4304 10013
rect 5172 10004 5224 10056
rect 7012 10072 7064 10124
rect 7748 10140 7800 10192
rect 8208 10208 8260 10260
rect 11520 10208 11572 10260
rect 12532 10208 12584 10260
rect 12992 10208 13044 10260
rect 13268 10208 13320 10260
rect 14188 10208 14240 10260
rect 15384 10208 15436 10260
rect 16120 10208 16172 10260
rect 15108 10140 15160 10192
rect 15844 10140 15896 10192
rect 16488 10208 16540 10260
rect 16764 10208 16816 10260
rect 16948 10208 17000 10260
rect 18420 10208 18472 10260
rect 1216 9868 1268 9920
rect 3516 9868 3568 9920
rect 4988 9936 5040 9988
rect 5356 9936 5408 9988
rect 5632 9936 5684 9988
rect 7104 9936 7156 9988
rect 7380 9936 7432 9988
rect 4712 9868 4764 9920
rect 4896 9868 4948 9920
rect 5724 9868 5776 9920
rect 6828 9868 6880 9920
rect 8944 10004 8996 10056
rect 9496 10072 9548 10124
rect 10048 10004 10100 10056
rect 15108 10004 15160 10056
rect 15292 10004 15344 10056
rect 16488 10004 16540 10056
rect 17684 10072 17736 10124
rect 7644 9868 7696 9920
rect 9496 9936 9548 9988
rect 13268 9936 13320 9988
rect 15384 9936 15436 9988
rect 17040 10047 17092 10056
rect 17040 10013 17049 10047
rect 17049 10013 17083 10047
rect 17083 10013 17092 10047
rect 17040 10004 17092 10013
rect 17500 10047 17552 10056
rect 17500 10013 17509 10047
rect 17509 10013 17543 10047
rect 17543 10013 17552 10047
rect 17500 10004 17552 10013
rect 16672 9936 16724 9988
rect 8944 9868 8996 9920
rect 12348 9868 12400 9920
rect 12624 9868 12676 9920
rect 12808 9868 12860 9920
rect 14832 9868 14884 9920
rect 17500 9868 17552 9920
rect 19064 10140 19116 10192
rect 18144 10072 18196 10124
rect 17776 9979 17828 9988
rect 17776 9945 17785 9979
rect 17785 9945 17819 9979
rect 17819 9945 17828 9979
rect 17776 9936 17828 9945
rect 18880 9936 18932 9988
rect 2610 9766 2662 9818
rect 2674 9766 2726 9818
rect 2738 9766 2790 9818
rect 2802 9766 2854 9818
rect 2866 9766 2918 9818
rect 7610 9766 7662 9818
rect 7674 9766 7726 9818
rect 7738 9766 7790 9818
rect 7802 9766 7854 9818
rect 7866 9766 7918 9818
rect 12610 9766 12662 9818
rect 12674 9766 12726 9818
rect 12738 9766 12790 9818
rect 12802 9766 12854 9818
rect 12866 9766 12918 9818
rect 17610 9766 17662 9818
rect 17674 9766 17726 9818
rect 17738 9766 17790 9818
rect 17802 9766 17854 9818
rect 17866 9766 17918 9818
rect 112 9664 164 9716
rect 1032 9596 1084 9648
rect 1584 9596 1636 9648
rect 2412 9664 2464 9716
rect 2596 9664 2648 9716
rect 388 9528 440 9580
rect 2872 9639 2924 9648
rect 2872 9605 2881 9639
rect 2881 9605 2915 9639
rect 2915 9605 2924 9639
rect 2872 9596 2924 9605
rect 2044 9571 2096 9580
rect 2044 9537 2053 9571
rect 2053 9537 2087 9571
rect 2087 9537 2096 9571
rect 2044 9528 2096 9537
rect 2412 9528 2464 9580
rect 2780 9528 2832 9580
rect 3792 9596 3844 9648
rect 4252 9664 4304 9716
rect 3056 9571 3108 9580
rect 3056 9537 3065 9571
rect 3065 9537 3099 9571
rect 3099 9537 3108 9571
rect 3056 9528 3108 9537
rect 2872 9460 2924 9512
rect 3884 9528 3936 9580
rect 3332 9503 3384 9512
rect 3332 9469 3341 9503
rect 3341 9469 3375 9503
rect 3375 9469 3384 9503
rect 3332 9460 3384 9469
rect 3516 9460 3568 9512
rect 4252 9460 4304 9512
rect 5632 9528 5684 9580
rect 5908 9664 5960 9716
rect 6184 9664 6236 9716
rect 6368 9664 6420 9716
rect 9036 9664 9088 9716
rect 10968 9664 11020 9716
rect 11060 9664 11112 9716
rect 12164 9664 12216 9716
rect 12256 9707 12308 9716
rect 12256 9673 12265 9707
rect 12265 9673 12299 9707
rect 12299 9673 12308 9707
rect 12256 9664 12308 9673
rect 13268 9664 13320 9716
rect 15108 9664 15160 9716
rect 17224 9664 17276 9716
rect 6828 9596 6880 9648
rect 6184 9528 6236 9580
rect 7104 9571 7156 9580
rect 7104 9537 7113 9571
rect 7113 9537 7147 9571
rect 7147 9537 7156 9571
rect 7104 9528 7156 9537
rect 5172 9460 5224 9512
rect 6368 9460 6420 9512
rect 7748 9571 7800 9580
rect 7748 9537 7757 9571
rect 7757 9537 7791 9571
rect 7791 9537 7800 9571
rect 7748 9528 7800 9537
rect 9036 9528 9088 9580
rect 9496 9528 9548 9580
rect 7656 9460 7708 9512
rect 7932 9460 7984 9512
rect 9772 9460 9824 9512
rect 10324 9571 10376 9580
rect 10324 9537 10333 9571
rect 10333 9537 10367 9571
rect 10367 9537 10376 9571
rect 10324 9528 10376 9537
rect 12348 9596 12400 9648
rect 12808 9596 12860 9648
rect 10600 9528 10652 9580
rect 10784 9528 10836 9580
rect 12532 9528 12584 9580
rect 14188 9571 14240 9586
rect 14188 9537 14197 9571
rect 14197 9537 14231 9571
rect 14231 9537 14240 9571
rect 14188 9534 14240 9537
rect 16948 9639 17000 9648
rect 16948 9605 16957 9639
rect 16957 9605 16991 9639
rect 16991 9605 17000 9639
rect 16948 9596 17000 9605
rect 2136 9392 2188 9444
rect 1676 9324 1728 9376
rect 2228 9324 2280 9376
rect 2688 9367 2740 9376
rect 2688 9333 2697 9367
rect 2697 9333 2731 9367
rect 2731 9333 2740 9367
rect 2688 9324 2740 9333
rect 3608 9324 3660 9376
rect 5172 9324 5224 9376
rect 6828 9324 6880 9376
rect 8208 9324 8260 9376
rect 9588 9392 9640 9444
rect 10876 9503 10928 9512
rect 10876 9469 10885 9503
rect 10885 9469 10919 9503
rect 10919 9469 10928 9503
rect 10876 9460 10928 9469
rect 11244 9460 11296 9512
rect 14464 9528 14516 9580
rect 14740 9528 14792 9580
rect 15108 9528 15160 9580
rect 15936 9528 15988 9580
rect 10968 9392 11020 9444
rect 12532 9392 12584 9444
rect 12992 9392 13044 9444
rect 15476 9460 15528 9512
rect 16212 9460 16264 9512
rect 16488 9528 16540 9580
rect 17408 9596 17460 9648
rect 17224 9571 17276 9580
rect 17224 9537 17233 9571
rect 17233 9537 17267 9571
rect 17267 9537 17276 9571
rect 17224 9528 17276 9537
rect 17776 9571 17828 9580
rect 17776 9537 17785 9571
rect 17785 9537 17819 9571
rect 17819 9537 17828 9571
rect 17776 9528 17828 9537
rect 18144 9571 18196 9580
rect 18144 9537 18153 9571
rect 18153 9537 18187 9571
rect 18187 9537 18196 9571
rect 18144 9528 18196 9537
rect 19340 9528 19392 9580
rect 14464 9435 14516 9444
rect 14464 9401 14473 9435
rect 14473 9401 14507 9435
rect 14507 9401 14516 9435
rect 14464 9392 14516 9401
rect 10600 9324 10652 9376
rect 10692 9324 10744 9376
rect 11704 9324 11756 9376
rect 11888 9324 11940 9376
rect 12348 9324 12400 9376
rect 14280 9324 14332 9376
rect 15936 9392 15988 9444
rect 14740 9324 14792 9376
rect 16488 9392 16540 9444
rect 16304 9324 16356 9376
rect 17776 9324 17828 9376
rect 1950 9222 2002 9274
rect 2014 9222 2066 9274
rect 2078 9222 2130 9274
rect 2142 9222 2194 9274
rect 2206 9222 2258 9274
rect 6950 9222 7002 9274
rect 7014 9222 7066 9274
rect 7078 9222 7130 9274
rect 7142 9222 7194 9274
rect 7206 9222 7258 9274
rect 11950 9222 12002 9274
rect 12014 9222 12066 9274
rect 12078 9222 12130 9274
rect 12142 9222 12194 9274
rect 12206 9222 12258 9274
rect 16950 9222 17002 9274
rect 17014 9222 17066 9274
rect 17078 9222 17130 9274
rect 17142 9222 17194 9274
rect 17206 9222 17258 9274
rect 2412 9120 2464 9172
rect 2504 9120 2556 9172
rect 3424 9120 3476 9172
rect 3792 9120 3844 9172
rect 4160 9120 4212 9172
rect 3884 9052 3936 9104
rect 5080 9120 5132 9172
rect 6828 9120 6880 9172
rect 7748 9120 7800 9172
rect 8392 9120 8444 9172
rect 9772 9120 9824 9172
rect 10692 9120 10744 9172
rect 11336 9120 11388 9172
rect 11612 9120 11664 9172
rect 12164 9120 12216 9172
rect 12440 9120 12492 9172
rect 13636 9120 13688 9172
rect 14464 9120 14516 9172
rect 10876 9052 10928 9104
rect 13728 9052 13780 9104
rect 13912 9052 13964 9104
rect 18236 9120 18288 9172
rect 14924 9052 14976 9104
rect 15200 9052 15252 9104
rect 1584 8959 1636 8968
rect 1584 8925 1593 8959
rect 1593 8925 1627 8959
rect 1627 8925 1636 8959
rect 1584 8916 1636 8925
rect 756 8848 808 8900
rect 1952 8959 2004 8968
rect 1952 8925 1961 8959
rect 1961 8925 1995 8959
rect 1995 8925 2004 8959
rect 1952 8916 2004 8925
rect 2964 8959 3016 8968
rect 2964 8925 2973 8959
rect 2973 8925 3007 8959
rect 3007 8925 3016 8959
rect 2964 8916 3016 8925
rect 7104 8984 7156 9036
rect 7380 8984 7432 9036
rect 2228 8891 2280 8900
rect 2228 8857 2237 8891
rect 2237 8857 2271 8891
rect 2271 8857 2280 8891
rect 2228 8848 2280 8857
rect 2412 8848 2464 8900
rect 4068 8916 4120 8968
rect 4160 8916 4212 8968
rect 4252 8916 4304 8968
rect 4620 8916 4672 8968
rect 3608 8848 3660 8900
rect 3884 8891 3936 8900
rect 3884 8857 3893 8891
rect 3893 8857 3927 8891
rect 3927 8857 3936 8891
rect 3884 8848 3936 8857
rect 5080 8959 5132 8968
rect 5080 8925 5089 8959
rect 5089 8925 5123 8959
rect 5123 8925 5132 8959
rect 5080 8916 5132 8925
rect 5264 8916 5316 8968
rect 5356 8916 5408 8968
rect 6368 8916 6420 8968
rect 8116 8984 8168 9036
rect 8576 8984 8628 9036
rect 9036 8984 9088 9036
rect 9220 8984 9272 9036
rect 7932 8848 7984 8900
rect 8116 8848 8168 8900
rect 9956 8848 10008 8900
rect 1124 8780 1176 8832
rect 1584 8780 1636 8832
rect 1860 8780 1912 8832
rect 2688 8780 2740 8832
rect 2780 8780 2832 8832
rect 4160 8780 4212 8832
rect 4252 8780 4304 8832
rect 4896 8780 4948 8832
rect 5356 8823 5408 8832
rect 5356 8789 5365 8823
rect 5365 8789 5399 8823
rect 5399 8789 5408 8823
rect 5356 8780 5408 8789
rect 7196 8780 7248 8832
rect 7840 8780 7892 8832
rect 8208 8780 8260 8832
rect 10324 8984 10376 9036
rect 11612 8984 11664 9036
rect 12624 8984 12676 9036
rect 16764 9052 16816 9104
rect 16396 8984 16448 9036
rect 17224 9052 17276 9104
rect 18696 9052 18748 9104
rect 10140 8916 10192 8968
rect 10324 8848 10376 8900
rect 12808 8916 12860 8968
rect 13636 8916 13688 8968
rect 14004 8916 14056 8968
rect 14188 8916 14240 8968
rect 16672 8916 16724 8968
rect 12532 8848 12584 8900
rect 16488 8848 16540 8900
rect 17224 8916 17276 8968
rect 10416 8823 10468 8832
rect 10416 8789 10425 8823
rect 10425 8789 10459 8823
rect 10459 8789 10468 8823
rect 10416 8780 10468 8789
rect 11888 8780 11940 8832
rect 12900 8780 12952 8832
rect 15108 8780 15160 8832
rect 16396 8780 16448 8832
rect 16764 8780 16816 8832
rect 17960 8780 18012 8832
rect 18420 8823 18472 8832
rect 18420 8789 18429 8823
rect 18429 8789 18463 8823
rect 18463 8789 18472 8823
rect 18420 8780 18472 8789
rect 2610 8678 2662 8730
rect 2674 8678 2726 8730
rect 2738 8678 2790 8730
rect 2802 8678 2854 8730
rect 2866 8678 2918 8730
rect 7610 8678 7662 8730
rect 7674 8678 7726 8730
rect 7738 8678 7790 8730
rect 7802 8678 7854 8730
rect 7866 8678 7918 8730
rect 12610 8678 12662 8730
rect 12674 8678 12726 8730
rect 12738 8678 12790 8730
rect 12802 8678 12854 8730
rect 12866 8678 12918 8730
rect 17610 8678 17662 8730
rect 17674 8678 17726 8730
rect 17738 8678 17790 8730
rect 17802 8678 17854 8730
rect 17866 8678 17918 8730
rect 1124 8576 1176 8628
rect 1676 8576 1728 8628
rect 2136 8619 2188 8628
rect 2136 8585 2145 8619
rect 2145 8585 2179 8619
rect 2179 8585 2188 8619
rect 2136 8576 2188 8585
rect 2228 8576 2280 8628
rect 2412 8576 2464 8628
rect 2596 8576 2648 8628
rect 1768 8508 1820 8560
rect 3884 8576 3936 8628
rect 4252 8576 4304 8628
rect 5264 8576 5316 8628
rect 6000 8576 6052 8628
rect 7104 8576 7156 8628
rect 7656 8576 7708 8628
rect 7748 8576 7800 8628
rect 8668 8576 8720 8628
rect 1676 8440 1728 8492
rect 204 8372 256 8424
rect 2412 8440 2464 8492
rect 3424 8508 3476 8560
rect 2320 8372 2372 8424
rect 2596 8415 2648 8424
rect 2596 8381 2605 8415
rect 2605 8381 2639 8415
rect 2639 8381 2648 8415
rect 2596 8372 2648 8381
rect 2964 8372 3016 8424
rect 3516 8440 3568 8492
rect 3884 8372 3936 8424
rect 4712 8508 4764 8560
rect 4252 8440 4304 8492
rect 5264 8372 5316 8424
rect 5724 8440 5776 8492
rect 6460 8440 6512 8492
rect 6552 8483 6604 8492
rect 6552 8449 6561 8483
rect 6561 8449 6595 8483
rect 6595 8449 6604 8483
rect 6552 8440 6604 8449
rect 6000 8415 6052 8424
rect 6000 8381 6009 8415
rect 6009 8381 6043 8415
rect 6043 8381 6052 8415
rect 6000 8372 6052 8381
rect 2228 8304 2280 8356
rect 2044 8236 2096 8288
rect 2320 8236 2372 8288
rect 4344 8304 4396 8356
rect 4804 8304 4856 8356
rect 6736 8483 6788 8492
rect 6736 8449 6745 8483
rect 6745 8449 6779 8483
rect 6779 8449 6788 8483
rect 6736 8440 6788 8449
rect 6828 8440 6880 8492
rect 7564 8440 7616 8492
rect 7656 8440 7708 8492
rect 8576 8440 8628 8492
rect 8668 8440 8720 8492
rect 9312 8483 9364 8492
rect 9312 8449 9321 8483
rect 9321 8449 9355 8483
rect 9355 8449 9364 8483
rect 9312 8440 9364 8449
rect 9588 8440 9640 8492
rect 10140 8576 10192 8628
rect 10692 8576 10744 8628
rect 13176 8576 13228 8628
rect 15108 8576 15160 8628
rect 16396 8576 16448 8628
rect 7840 8372 7892 8424
rect 9772 8372 9824 8424
rect 8576 8304 8628 8356
rect 10324 8483 10376 8492
rect 10324 8449 10333 8483
rect 10333 8449 10367 8483
rect 10367 8449 10376 8483
rect 10324 8440 10376 8449
rect 11336 8508 11388 8560
rect 12164 8508 12216 8560
rect 13728 8508 13780 8560
rect 14004 8508 14056 8560
rect 15752 8508 15804 8560
rect 10968 8440 11020 8492
rect 12256 8440 12308 8492
rect 15384 8440 15436 8492
rect 18788 8508 18840 8560
rect 18052 8440 18104 8492
rect 10232 8372 10284 8424
rect 15476 8372 15528 8424
rect 15660 8372 15712 8424
rect 19524 8372 19576 8424
rect 10416 8304 10468 8356
rect 10600 8347 10652 8356
rect 10600 8313 10609 8347
rect 10609 8313 10643 8347
rect 10643 8313 10652 8347
rect 10600 8304 10652 8313
rect 11336 8304 11388 8356
rect 2688 8236 2740 8288
rect 3056 8236 3108 8288
rect 5080 8236 5132 8288
rect 5540 8236 5592 8288
rect 7012 8236 7064 8288
rect 8116 8236 8168 8288
rect 8760 8236 8812 8288
rect 9312 8236 9364 8288
rect 9404 8236 9456 8288
rect 9680 8236 9732 8288
rect 9956 8236 10008 8288
rect 10692 8236 10744 8288
rect 11152 8236 11204 8288
rect 12808 8236 12860 8288
rect 13728 8304 13780 8356
rect 14556 8304 14608 8356
rect 14924 8236 14976 8288
rect 15476 8236 15528 8288
rect 17592 8236 17644 8288
rect 1950 8134 2002 8186
rect 2014 8134 2066 8186
rect 2078 8134 2130 8186
rect 2142 8134 2194 8186
rect 2206 8134 2258 8186
rect 6950 8134 7002 8186
rect 7014 8134 7066 8186
rect 7078 8134 7130 8186
rect 7142 8134 7194 8186
rect 7206 8134 7258 8186
rect 11950 8134 12002 8186
rect 12014 8134 12066 8186
rect 12078 8134 12130 8186
rect 12142 8134 12194 8186
rect 12206 8134 12258 8186
rect 16950 8134 17002 8186
rect 17014 8134 17066 8186
rect 17078 8134 17130 8186
rect 17142 8134 17194 8186
rect 17206 8134 17258 8186
rect 2780 8032 2832 8084
rect 4620 8032 4672 8084
rect 5264 8032 5316 8084
rect 756 7964 808 8016
rect 2872 7964 2924 8016
rect 6276 7964 6328 8016
rect 3608 7896 3660 7948
rect 3884 7896 3936 7948
rect 12440 8032 12492 8084
rect 13912 8032 13964 8084
rect 16028 8032 16080 8084
rect 1768 7760 1820 7812
rect 3884 7760 3936 7812
rect 4344 7803 4396 7812
rect 4344 7769 4353 7803
rect 4353 7769 4387 7803
rect 4387 7769 4396 7803
rect 4344 7760 4396 7769
rect 1308 7692 1360 7744
rect 2780 7692 2832 7744
rect 3056 7692 3108 7744
rect 4528 7871 4580 7880
rect 4528 7837 4537 7871
rect 4537 7837 4571 7871
rect 4571 7837 4580 7871
rect 4528 7828 4580 7837
rect 6000 7871 6052 7880
rect 6000 7837 6009 7871
rect 6009 7837 6043 7871
rect 6043 7837 6052 7871
rect 6644 7896 6696 7948
rect 6000 7828 6052 7837
rect 6736 7871 6788 7880
rect 6736 7837 6745 7871
rect 6745 7837 6779 7871
rect 6779 7837 6788 7871
rect 6736 7828 6788 7837
rect 7196 7939 7248 7948
rect 7196 7905 7205 7939
rect 7205 7905 7239 7939
rect 7239 7905 7248 7939
rect 7196 7896 7248 7905
rect 7288 7896 7340 7948
rect 7932 7896 7984 7948
rect 11244 7964 11296 8016
rect 13360 7964 13412 8016
rect 15108 7964 15160 8016
rect 9956 7896 10008 7948
rect 10692 7896 10744 7948
rect 12992 7896 13044 7948
rect 7564 7828 7616 7880
rect 7840 7828 7892 7880
rect 8208 7828 8260 7880
rect 8392 7828 8444 7880
rect 7012 7692 7064 7744
rect 7196 7760 7248 7812
rect 9128 7828 9180 7880
rect 9312 7871 9364 7880
rect 9312 7837 9321 7871
rect 9321 7837 9355 7871
rect 9355 7837 9364 7871
rect 9312 7828 9364 7837
rect 9772 7871 9824 7880
rect 9772 7837 9781 7871
rect 9781 7837 9815 7871
rect 9815 7837 9824 7871
rect 9772 7828 9824 7837
rect 10784 7828 10836 7880
rect 8116 7692 8168 7744
rect 13820 7828 13872 7880
rect 13912 7828 13964 7880
rect 14832 7828 14884 7880
rect 13728 7760 13780 7812
rect 10784 7692 10836 7744
rect 11152 7692 11204 7744
rect 11520 7692 11572 7744
rect 12624 7692 12676 7744
rect 12808 7692 12860 7744
rect 13360 7692 13412 7744
rect 15384 7871 15436 7880
rect 15384 7837 15393 7871
rect 15393 7837 15427 7871
rect 15427 7837 15436 7871
rect 15384 7828 15436 7837
rect 15476 7871 15528 7880
rect 15476 7837 15485 7871
rect 15485 7837 15519 7871
rect 15519 7837 15528 7871
rect 15476 7828 15528 7837
rect 15844 7964 15896 8016
rect 16764 8032 16816 8084
rect 16212 7896 16264 7948
rect 16120 7871 16172 7880
rect 16120 7837 16129 7871
rect 16129 7837 16163 7871
rect 16163 7837 16172 7871
rect 16120 7828 16172 7837
rect 17040 7828 17092 7880
rect 18144 7828 18196 7880
rect 17224 7760 17276 7812
rect 19064 7760 19116 7812
rect 15844 7692 15896 7744
rect 16304 7735 16356 7744
rect 16304 7701 16313 7735
rect 16313 7701 16347 7735
rect 16347 7701 16356 7735
rect 16304 7692 16356 7701
rect 2610 7590 2662 7642
rect 2674 7590 2726 7642
rect 2738 7590 2790 7642
rect 2802 7590 2854 7642
rect 2866 7590 2918 7642
rect 7610 7590 7662 7642
rect 7674 7590 7726 7642
rect 7738 7590 7790 7642
rect 7802 7590 7854 7642
rect 7866 7590 7918 7642
rect 12610 7590 12662 7642
rect 12674 7590 12726 7642
rect 12738 7590 12790 7642
rect 12802 7590 12854 7642
rect 12866 7590 12918 7642
rect 17610 7590 17662 7642
rect 17674 7590 17726 7642
rect 17738 7590 17790 7642
rect 17802 7590 17854 7642
rect 17866 7590 17918 7642
rect 4712 7488 4764 7540
rect 5264 7488 5316 7540
rect 8392 7488 8444 7540
rect 8852 7488 8904 7540
rect 9588 7488 9640 7540
rect 9772 7488 9824 7540
rect 10600 7488 10652 7540
rect 10876 7488 10928 7540
rect 11520 7488 11572 7540
rect 13084 7488 13136 7540
rect 1492 7420 1544 7472
rect 4896 7420 4948 7472
rect 6276 7420 6328 7472
rect 4344 7352 4396 7404
rect 7564 7395 7616 7404
rect 7564 7361 7573 7395
rect 7573 7361 7607 7395
rect 7607 7361 7616 7395
rect 7564 7352 7616 7361
rect 8300 7420 8352 7472
rect 4528 7327 4580 7336
rect 4528 7293 4537 7327
rect 4537 7293 4571 7327
rect 4571 7293 4580 7327
rect 4528 7284 4580 7293
rect 6276 7284 6328 7336
rect 6920 7284 6972 7336
rect 7104 7284 7156 7336
rect 7656 7284 7708 7336
rect 8116 7352 8168 7404
rect 8668 7352 8720 7404
rect 11060 7420 11112 7472
rect 16304 7488 16356 7540
rect 15108 7420 15160 7472
rect 17224 7420 17276 7472
rect 9680 7352 9732 7404
rect 9864 7395 9916 7404
rect 9864 7361 9873 7395
rect 9873 7361 9907 7395
rect 9907 7361 9916 7395
rect 9864 7352 9916 7361
rect 10232 7352 10284 7404
rect 8852 7284 8904 7336
rect 9956 7327 10008 7336
rect 9956 7293 9965 7327
rect 9965 7293 9999 7327
rect 9999 7293 10008 7327
rect 9956 7284 10008 7293
rect 2504 7216 2556 7268
rect 5540 7216 5592 7268
rect 7012 7216 7064 7268
rect 10784 7352 10836 7404
rect 11520 7395 11572 7404
rect 11520 7361 11529 7395
rect 11529 7361 11563 7395
rect 11563 7361 11572 7395
rect 11520 7352 11572 7361
rect 11612 7352 11664 7404
rect 11980 7352 12032 7404
rect 14372 7395 14424 7404
rect 14372 7361 14381 7395
rect 14381 7361 14415 7395
rect 14415 7361 14424 7395
rect 14372 7352 14424 7361
rect 14464 7352 14516 7404
rect 17040 7395 17092 7404
rect 17040 7361 17049 7395
rect 17049 7361 17083 7395
rect 17083 7361 17092 7395
rect 17040 7352 17092 7361
rect 10600 7284 10652 7336
rect 12348 7284 12400 7336
rect 15752 7284 15804 7336
rect 3976 7148 4028 7200
rect 8392 7148 8444 7200
rect 12992 7216 13044 7268
rect 13728 7216 13780 7268
rect 13912 7216 13964 7268
rect 17960 7216 18012 7268
rect 10600 7148 10652 7200
rect 11152 7148 11204 7200
rect 11336 7148 11388 7200
rect 12256 7148 12308 7200
rect 1950 7046 2002 7098
rect 2014 7046 2066 7098
rect 2078 7046 2130 7098
rect 2142 7046 2194 7098
rect 2206 7046 2258 7098
rect 6950 7046 7002 7098
rect 7014 7046 7066 7098
rect 7078 7046 7130 7098
rect 7142 7046 7194 7098
rect 7206 7046 7258 7098
rect 11950 7046 12002 7098
rect 12014 7046 12066 7098
rect 12078 7046 12130 7098
rect 12142 7046 12194 7098
rect 12206 7046 12258 7098
rect 16950 7046 17002 7098
rect 17014 7046 17066 7098
rect 17078 7046 17130 7098
rect 17142 7046 17194 7098
rect 17206 7046 17258 7098
rect 112 6944 164 6996
rect 1768 6944 1820 6996
rect 2504 6944 2556 6996
rect 3148 6944 3200 6996
rect 3424 6944 3476 6996
rect 4068 6944 4120 6996
rect 4344 6944 4396 6996
rect 3884 6876 3936 6928
rect 2320 6808 2372 6860
rect 3608 6808 3660 6860
rect 4344 6808 4396 6860
rect 5724 6944 5776 6996
rect 8024 6944 8076 6996
rect 8116 6944 8168 6996
rect 8760 6944 8812 6996
rect 5816 6876 5868 6928
rect 6460 6876 6512 6928
rect 8300 6876 8352 6928
rect 8392 6876 8444 6928
rect 15844 6944 15896 6996
rect 8944 6876 8996 6928
rect 6092 6808 6144 6860
rect 1492 6715 1544 6724
rect 1492 6681 1501 6715
rect 1501 6681 1535 6715
rect 1535 6681 1544 6715
rect 1492 6672 1544 6681
rect 3148 6672 3200 6724
rect 3332 6672 3384 6724
rect 3792 6740 3844 6792
rect 4068 6783 4120 6792
rect 4068 6749 4077 6783
rect 4077 6749 4111 6783
rect 4111 6749 4120 6783
rect 4068 6740 4120 6749
rect 4436 6783 4488 6792
rect 4436 6749 4445 6783
rect 4445 6749 4479 6783
rect 4479 6749 4488 6783
rect 4436 6740 4488 6749
rect 6644 6783 6696 6792
rect 6644 6749 6653 6783
rect 6653 6749 6687 6783
rect 6687 6749 6696 6783
rect 6644 6740 6696 6749
rect 7564 6740 7616 6792
rect 7656 6783 7708 6792
rect 7656 6749 7665 6783
rect 7665 6749 7699 6783
rect 7699 6749 7708 6783
rect 7656 6740 7708 6749
rect 8024 6783 8076 6792
rect 4804 6672 4856 6724
rect 5816 6672 5868 6724
rect 3792 6604 3844 6656
rect 5080 6604 5132 6656
rect 7196 6604 7248 6656
rect 8024 6749 8033 6783
rect 8033 6749 8067 6783
rect 8067 6749 8076 6783
rect 8024 6740 8076 6749
rect 8116 6783 8168 6792
rect 8116 6749 8125 6783
rect 8125 6749 8159 6783
rect 8159 6749 8168 6783
rect 8116 6740 8168 6749
rect 8208 6783 8260 6792
rect 8208 6749 8217 6783
rect 8217 6749 8251 6783
rect 8251 6749 8260 6783
rect 8208 6740 8260 6749
rect 8852 6808 8904 6860
rect 9496 6808 9548 6860
rect 12808 6808 12860 6860
rect 8392 6783 8444 6792
rect 8392 6749 8401 6783
rect 8401 6749 8435 6783
rect 8435 6749 8444 6783
rect 8392 6740 8444 6749
rect 10876 6740 10928 6792
rect 11060 6740 11112 6792
rect 11612 6740 11664 6792
rect 12532 6740 12584 6792
rect 12624 6783 12676 6792
rect 12624 6749 12633 6783
rect 12633 6749 12667 6783
rect 12667 6749 12676 6783
rect 12624 6740 12676 6749
rect 13544 6876 13596 6928
rect 14832 6876 14884 6928
rect 12992 6808 13044 6860
rect 19248 6808 19300 6860
rect 17500 6740 17552 6792
rect 19432 6740 19484 6792
rect 12256 6672 12308 6724
rect 7932 6604 7984 6656
rect 8208 6604 8260 6656
rect 8300 6604 8352 6656
rect 8760 6604 8812 6656
rect 9680 6604 9732 6656
rect 10784 6604 10836 6656
rect 12532 6604 12584 6656
rect 12808 6604 12860 6656
rect 16856 6672 16908 6724
rect 14004 6604 14056 6656
rect 14740 6604 14792 6656
rect 18420 6647 18472 6656
rect 18420 6613 18429 6647
rect 18429 6613 18463 6647
rect 18463 6613 18472 6647
rect 18420 6604 18472 6613
rect 2610 6502 2662 6554
rect 2674 6502 2726 6554
rect 2738 6502 2790 6554
rect 2802 6502 2854 6554
rect 2866 6502 2918 6554
rect 7610 6502 7662 6554
rect 7674 6502 7726 6554
rect 7738 6502 7790 6554
rect 7802 6502 7854 6554
rect 7866 6502 7918 6554
rect 12610 6502 12662 6554
rect 12674 6502 12726 6554
rect 12738 6502 12790 6554
rect 12802 6502 12854 6554
rect 12866 6502 12918 6554
rect 17610 6502 17662 6554
rect 17674 6502 17726 6554
rect 17738 6502 17790 6554
rect 17802 6502 17854 6554
rect 17866 6502 17918 6554
rect 4252 6443 4304 6452
rect 4252 6409 4279 6443
rect 4279 6409 4304 6443
rect 4252 6400 4304 6409
rect 5540 6400 5592 6452
rect 7564 6400 7616 6452
rect 2872 6332 2924 6384
rect 3148 6332 3200 6384
rect 3332 6332 3384 6384
rect 3516 6332 3568 6384
rect 3608 6307 3660 6316
rect 3608 6273 3617 6307
rect 3617 6273 3651 6307
rect 3651 6273 3660 6307
rect 3608 6264 3660 6273
rect 3148 6196 3200 6248
rect 3976 6307 4028 6316
rect 3976 6273 3985 6307
rect 3985 6273 4019 6307
rect 4019 6273 4028 6307
rect 3976 6264 4028 6273
rect 572 6128 624 6180
rect 2596 6128 2648 6180
rect 1584 6060 1636 6112
rect 3976 6128 4028 6180
rect 4436 6375 4488 6384
rect 4436 6341 4445 6375
rect 4445 6341 4479 6375
rect 4479 6341 4488 6375
rect 4436 6332 4488 6341
rect 4896 6332 4948 6384
rect 7656 6332 7708 6384
rect 7932 6400 7984 6452
rect 8116 6400 8168 6452
rect 8576 6400 8628 6452
rect 9680 6400 9732 6452
rect 11704 6400 11756 6452
rect 14096 6400 14148 6452
rect 15936 6400 15988 6452
rect 17592 6400 17644 6452
rect 4436 6196 4488 6248
rect 5080 6264 5132 6316
rect 5724 6307 5776 6316
rect 5724 6273 5733 6307
rect 5733 6273 5767 6307
rect 5767 6273 5776 6307
rect 5724 6264 5776 6273
rect 6184 6264 6236 6316
rect 6644 6264 6696 6316
rect 7288 6264 7340 6316
rect 10048 6332 10100 6384
rect 10232 6375 10284 6384
rect 10232 6341 10241 6375
rect 10241 6341 10275 6375
rect 10275 6341 10284 6375
rect 10232 6332 10284 6341
rect 10968 6332 11020 6384
rect 11796 6332 11848 6384
rect 8116 6307 8168 6316
rect 8116 6273 8125 6307
rect 8125 6273 8159 6307
rect 8159 6273 8168 6307
rect 8116 6264 8168 6273
rect 8208 6264 8260 6316
rect 7104 6196 7156 6248
rect 7564 6196 7616 6248
rect 5540 6128 5592 6180
rect 8116 6128 8168 6180
rect 9496 6239 9548 6248
rect 9496 6205 9505 6239
rect 9505 6205 9539 6239
rect 9539 6205 9548 6239
rect 9496 6196 9548 6205
rect 9680 6307 9732 6316
rect 9680 6273 9689 6307
rect 9689 6273 9723 6307
rect 9723 6273 9732 6307
rect 9680 6264 9732 6273
rect 10692 6264 10744 6316
rect 10784 6264 10836 6316
rect 15476 6332 15528 6384
rect 12256 6264 12308 6316
rect 13360 6264 13412 6316
rect 17960 6264 18012 6316
rect 12440 6196 12492 6248
rect 14648 6196 14700 6248
rect 14924 6128 14976 6180
rect 15752 6128 15804 6180
rect 3516 6060 3568 6112
rect 4620 6060 4672 6112
rect 4988 6060 5040 6112
rect 6276 6060 6328 6112
rect 7656 6060 7708 6112
rect 8944 6060 8996 6112
rect 11244 6060 11296 6112
rect 14464 6060 14516 6112
rect 14648 6060 14700 6112
rect 16580 6060 16632 6112
rect 1950 5958 2002 6010
rect 2014 5958 2066 6010
rect 2078 5958 2130 6010
rect 2142 5958 2194 6010
rect 2206 5958 2258 6010
rect 6950 5958 7002 6010
rect 7014 5958 7066 6010
rect 7078 5958 7130 6010
rect 7142 5958 7194 6010
rect 7206 5958 7258 6010
rect 11950 5958 12002 6010
rect 12014 5958 12066 6010
rect 12078 5958 12130 6010
rect 12142 5958 12194 6010
rect 12206 5958 12258 6010
rect 16950 5958 17002 6010
rect 17014 5958 17066 6010
rect 17078 5958 17130 6010
rect 17142 5958 17194 6010
rect 17206 5958 17258 6010
rect 2504 5856 2556 5908
rect 2688 5856 2740 5908
rect 3332 5856 3384 5908
rect 3608 5856 3660 5908
rect 1400 5788 1452 5840
rect 7840 5856 7892 5908
rect 8852 5856 8904 5908
rect 8944 5899 8996 5908
rect 8944 5865 8953 5899
rect 8953 5865 8987 5899
rect 8987 5865 8996 5899
rect 8944 5856 8996 5865
rect 10140 5856 10192 5908
rect 10508 5899 10560 5908
rect 10508 5865 10517 5899
rect 10517 5865 10551 5899
rect 10551 5865 10560 5899
rect 10508 5856 10560 5865
rect 10876 5856 10928 5908
rect 12624 5856 12676 5908
rect 9128 5788 9180 5840
rect 848 5720 900 5772
rect 2872 5720 2924 5772
rect 2412 5695 2464 5704
rect 2412 5661 2421 5695
rect 2421 5661 2455 5695
rect 2455 5661 2464 5695
rect 2412 5652 2464 5661
rect 2596 5652 2648 5704
rect 756 5584 808 5636
rect 1308 5516 1360 5568
rect 1492 5516 1544 5568
rect 2320 5584 2372 5636
rect 3424 5720 3476 5772
rect 4068 5720 4120 5772
rect 4804 5720 4856 5772
rect 4896 5720 4948 5772
rect 6000 5720 6052 5772
rect 6644 5763 6696 5772
rect 6644 5729 6653 5763
rect 6653 5729 6687 5763
rect 6687 5729 6696 5763
rect 6644 5720 6696 5729
rect 6828 5720 6880 5772
rect 4528 5652 4580 5704
rect 6460 5652 6512 5704
rect 7472 5695 7524 5704
rect 7472 5661 7481 5695
rect 7481 5661 7515 5695
rect 7515 5661 7524 5695
rect 7472 5652 7524 5661
rect 7656 5652 7708 5704
rect 8300 5652 8352 5704
rect 8944 5652 8996 5704
rect 9128 5695 9180 5704
rect 9128 5661 9137 5695
rect 9137 5661 9171 5695
rect 9171 5661 9180 5695
rect 9128 5652 9180 5661
rect 3608 5516 3660 5568
rect 4160 5516 4212 5568
rect 5264 5516 5316 5568
rect 5816 5516 5868 5568
rect 6736 5516 6788 5568
rect 7840 5516 7892 5568
rect 7932 5516 7984 5568
rect 8208 5516 8260 5568
rect 8392 5584 8444 5636
rect 13544 5720 13596 5772
rect 9956 5652 10008 5704
rect 10600 5652 10652 5704
rect 9772 5584 9824 5636
rect 11152 5652 11204 5704
rect 11704 5652 11756 5704
rect 11796 5695 11848 5704
rect 11796 5661 11805 5695
rect 11805 5661 11839 5695
rect 11839 5661 11848 5695
rect 11796 5652 11848 5661
rect 13176 5652 13228 5704
rect 14004 5720 14056 5772
rect 15108 5788 15160 5840
rect 16856 5856 16908 5908
rect 16028 5788 16080 5840
rect 14464 5763 14516 5772
rect 14464 5729 14473 5763
rect 14473 5729 14507 5763
rect 14507 5729 14516 5763
rect 14464 5720 14516 5729
rect 14832 5763 14884 5772
rect 14832 5729 14841 5763
rect 14841 5729 14875 5763
rect 14875 5729 14884 5763
rect 14832 5720 14884 5729
rect 16488 5720 16540 5772
rect 16580 5763 16632 5772
rect 16580 5729 16589 5763
rect 16589 5729 16623 5763
rect 16623 5729 16632 5763
rect 16580 5720 16632 5729
rect 15108 5652 15160 5704
rect 15200 5695 15252 5704
rect 15200 5661 15209 5695
rect 15209 5661 15243 5695
rect 15243 5661 15252 5695
rect 15200 5652 15252 5661
rect 9128 5516 9180 5568
rect 10600 5516 10652 5568
rect 10784 5516 10836 5568
rect 11612 5516 11664 5568
rect 14188 5559 14240 5568
rect 14188 5525 14197 5559
rect 14197 5525 14231 5559
rect 14231 5525 14240 5559
rect 14188 5516 14240 5525
rect 14924 5584 14976 5636
rect 16304 5652 16356 5704
rect 16764 5695 16816 5704
rect 16764 5661 16773 5695
rect 16773 5661 16807 5695
rect 16807 5661 16816 5695
rect 16764 5652 16816 5661
rect 16580 5584 16632 5636
rect 14832 5516 14884 5568
rect 15200 5516 15252 5568
rect 17960 5856 18012 5908
rect 17316 5720 17368 5772
rect 17592 5695 17644 5704
rect 17592 5661 17601 5695
rect 17601 5661 17635 5695
rect 17635 5661 17644 5695
rect 17592 5652 17644 5661
rect 18328 5584 18380 5636
rect 2610 5414 2662 5466
rect 2674 5414 2726 5466
rect 2738 5414 2790 5466
rect 2802 5414 2854 5466
rect 2866 5414 2918 5466
rect 7610 5414 7662 5466
rect 7674 5414 7726 5466
rect 7738 5414 7790 5466
rect 7802 5414 7854 5466
rect 7866 5414 7918 5466
rect 12610 5414 12662 5466
rect 12674 5414 12726 5466
rect 12738 5414 12790 5466
rect 12802 5414 12854 5466
rect 12866 5414 12918 5466
rect 17610 5414 17662 5466
rect 17674 5414 17726 5466
rect 17738 5414 17790 5466
rect 17802 5414 17854 5466
rect 17866 5414 17918 5466
rect 1124 5312 1176 5364
rect 1308 5312 1360 5364
rect 3056 5312 3108 5364
rect 2412 5244 2464 5296
rect 3424 5244 3476 5296
rect 3608 5244 3660 5296
rect 3056 5176 3108 5228
rect 3976 5176 4028 5228
rect 4160 5219 4212 5228
rect 4160 5185 4169 5219
rect 4169 5185 4203 5219
rect 4203 5185 4212 5219
rect 4160 5176 4212 5185
rect 4344 5176 4396 5228
rect 4068 5151 4120 5160
rect 4068 5117 4077 5151
rect 4077 5117 4111 5151
rect 4111 5117 4120 5151
rect 4068 5108 4120 5117
rect 5908 5244 5960 5296
rect 4988 5219 5040 5228
rect 4988 5185 4997 5219
rect 4997 5185 5031 5219
rect 5031 5185 5040 5219
rect 4988 5176 5040 5185
rect 5172 5219 5224 5228
rect 5172 5185 5181 5219
rect 5181 5185 5215 5219
rect 5215 5185 5224 5219
rect 5172 5176 5224 5185
rect 5632 5219 5684 5228
rect 5632 5185 5641 5219
rect 5641 5185 5675 5219
rect 5675 5185 5684 5219
rect 5632 5176 5684 5185
rect 7288 5355 7340 5364
rect 7288 5321 7297 5355
rect 7297 5321 7331 5355
rect 7331 5321 7340 5355
rect 7288 5312 7340 5321
rect 7472 5312 7524 5364
rect 7748 5312 7800 5364
rect 10600 5312 10652 5364
rect 10876 5312 10928 5364
rect 11520 5312 11572 5364
rect 6460 5176 6512 5228
rect 4160 5040 4212 5092
rect 4804 5083 4856 5092
rect 4804 5049 4813 5083
rect 4813 5049 4847 5083
rect 4847 5049 4856 5083
rect 4804 5040 4856 5049
rect 4344 4972 4396 5024
rect 5264 5040 5316 5092
rect 7288 5176 7340 5228
rect 7932 5219 7984 5228
rect 7932 5185 7941 5219
rect 7941 5185 7975 5219
rect 7975 5185 7984 5219
rect 7932 5176 7984 5185
rect 8116 5176 8168 5228
rect 8852 5287 8904 5296
rect 8852 5253 8861 5287
rect 8861 5253 8895 5287
rect 8895 5253 8904 5287
rect 8852 5244 8904 5253
rect 10416 5244 10468 5296
rect 10508 5244 10560 5296
rect 9036 5219 9088 5228
rect 9036 5185 9045 5219
rect 9045 5185 9079 5219
rect 9079 5185 9088 5219
rect 9036 5176 9088 5185
rect 9128 5176 9180 5228
rect 10968 5176 11020 5228
rect 12532 5244 12584 5296
rect 16396 5312 16448 5364
rect 16488 5244 16540 5296
rect 17500 5355 17552 5364
rect 17500 5321 17509 5355
rect 17509 5321 17543 5355
rect 17543 5321 17552 5355
rect 17500 5312 17552 5321
rect 12256 5176 12308 5228
rect 13452 5176 13504 5228
rect 15476 5219 15528 5228
rect 15476 5185 15485 5219
rect 15485 5185 15519 5219
rect 15519 5185 15528 5219
rect 15476 5176 15528 5185
rect 15660 5219 15712 5228
rect 15660 5185 15669 5219
rect 15669 5185 15703 5219
rect 15703 5185 15712 5219
rect 15660 5176 15712 5185
rect 7012 5151 7064 5160
rect 7012 5117 7021 5151
rect 7021 5117 7055 5151
rect 7055 5117 7064 5151
rect 7012 5108 7064 5117
rect 7472 5108 7524 5160
rect 8944 5108 8996 5160
rect 5724 5015 5776 5024
rect 5724 4981 5733 5015
rect 5733 4981 5767 5015
rect 5767 4981 5776 5015
rect 5724 4972 5776 4981
rect 6000 4972 6052 5024
rect 6736 4972 6788 5024
rect 8392 5040 8444 5092
rect 8668 5040 8720 5092
rect 8300 4972 8352 5024
rect 11796 5108 11848 5160
rect 13084 5108 13136 5160
rect 16120 5108 16172 5160
rect 16488 5151 16540 5160
rect 16488 5117 16497 5151
rect 16497 5117 16531 5151
rect 16531 5117 16540 5151
rect 16488 5108 16540 5117
rect 16672 5108 16724 5160
rect 16764 5108 16816 5160
rect 17960 5176 18012 5228
rect 18328 5219 18380 5228
rect 18328 5185 18337 5219
rect 18337 5185 18371 5219
rect 18371 5185 18380 5219
rect 18328 5176 18380 5185
rect 10048 5040 10100 5092
rect 10600 4972 10652 5024
rect 12256 4972 12308 5024
rect 12532 4972 12584 5024
rect 16672 4972 16724 5024
rect 18328 5015 18380 5024
rect 18328 4981 18337 5015
rect 18337 4981 18371 5015
rect 18371 4981 18380 5015
rect 18328 4972 18380 4981
rect 1950 4870 2002 4922
rect 2014 4870 2066 4922
rect 2078 4870 2130 4922
rect 2142 4870 2194 4922
rect 2206 4870 2258 4922
rect 6950 4870 7002 4922
rect 7014 4870 7066 4922
rect 7078 4870 7130 4922
rect 7142 4870 7194 4922
rect 7206 4870 7258 4922
rect 11950 4870 12002 4922
rect 12014 4870 12066 4922
rect 12078 4870 12130 4922
rect 12142 4870 12194 4922
rect 12206 4870 12258 4922
rect 16950 4870 17002 4922
rect 17014 4870 17066 4922
rect 17078 4870 17130 4922
rect 17142 4870 17194 4922
rect 17206 4870 17258 4922
rect 1768 4768 1820 4820
rect 1952 4768 2004 4820
rect 2504 4768 2556 4820
rect 5080 4768 5132 4820
rect 5448 4768 5500 4820
rect 5816 4768 5868 4820
rect 6736 4768 6788 4820
rect 2780 4743 2832 4752
rect 2780 4709 2789 4743
rect 2789 4709 2823 4743
rect 2823 4709 2832 4743
rect 2780 4700 2832 4709
rect 1768 4632 1820 4684
rect 2412 4564 2464 4616
rect 4252 4700 4304 4752
rect 5172 4700 5224 4752
rect 3240 4632 3292 4684
rect 4436 4632 4488 4684
rect 4712 4632 4764 4684
rect 7012 4700 7064 4752
rect 7380 4768 7432 4820
rect 9956 4768 10008 4820
rect 12072 4768 12124 4820
rect 7196 4700 7248 4752
rect 9128 4700 9180 4752
rect 9680 4700 9732 4752
rect 14648 4811 14700 4820
rect 14648 4777 14657 4811
rect 14657 4777 14691 4811
rect 14691 4777 14700 4811
rect 14648 4768 14700 4777
rect 15292 4768 15344 4820
rect 14832 4700 14884 4752
rect 3976 4607 4028 4616
rect 3976 4573 3985 4607
rect 3985 4573 4019 4607
rect 4019 4573 4028 4607
rect 3976 4564 4028 4573
rect 4160 4564 4212 4616
rect 4344 4496 4396 4548
rect 4712 4496 4764 4548
rect 5540 4607 5592 4616
rect 5540 4573 5549 4607
rect 5549 4573 5583 4607
rect 5583 4573 5592 4607
rect 5540 4564 5592 4573
rect 6092 4428 6144 4480
rect 7196 4607 7248 4616
rect 7196 4573 7205 4607
rect 7205 4573 7239 4607
rect 7239 4573 7248 4607
rect 7196 4564 7248 4573
rect 6828 4496 6880 4548
rect 7748 4564 7800 4616
rect 8024 4564 8076 4616
rect 8116 4564 8168 4616
rect 8576 4564 8628 4616
rect 10416 4607 10468 4616
rect 10416 4573 10425 4607
rect 10425 4573 10459 4607
rect 10459 4573 10468 4607
rect 10416 4564 10468 4573
rect 10692 4564 10744 4616
rect 11520 4607 11572 4616
rect 11520 4573 11529 4607
rect 11529 4573 11563 4607
rect 11563 4573 11572 4607
rect 11520 4564 11572 4573
rect 11796 4607 11848 4616
rect 11796 4573 11805 4607
rect 11805 4573 11839 4607
rect 11839 4573 11848 4607
rect 11796 4564 11848 4573
rect 11888 4564 11940 4616
rect 13544 4564 13596 4616
rect 8852 4496 8904 4548
rect 9956 4496 10008 4548
rect 13268 4496 13320 4548
rect 14556 4607 14608 4616
rect 14556 4573 14565 4607
rect 14565 4573 14599 4607
rect 14599 4573 14608 4607
rect 14556 4564 14608 4573
rect 14648 4607 14700 4616
rect 14648 4573 14657 4607
rect 14657 4573 14691 4607
rect 14691 4573 14700 4607
rect 14648 4564 14700 4573
rect 14740 4564 14792 4616
rect 15016 4607 15068 4616
rect 15016 4573 15025 4607
rect 15025 4573 15059 4607
rect 15059 4573 15068 4607
rect 15016 4564 15068 4573
rect 15936 4632 15988 4684
rect 16120 4564 16172 4616
rect 16304 4564 16356 4616
rect 8760 4428 8812 4480
rect 10692 4428 10744 4480
rect 18972 4428 19024 4480
rect 2610 4326 2662 4378
rect 2674 4326 2726 4378
rect 2738 4326 2790 4378
rect 2802 4326 2854 4378
rect 2866 4326 2918 4378
rect 7610 4326 7662 4378
rect 7674 4326 7726 4378
rect 7738 4326 7790 4378
rect 7802 4326 7854 4378
rect 7866 4326 7918 4378
rect 12610 4326 12662 4378
rect 12674 4326 12726 4378
rect 12738 4326 12790 4378
rect 12802 4326 12854 4378
rect 12866 4326 12918 4378
rect 17610 4326 17662 4378
rect 17674 4326 17726 4378
rect 17738 4326 17790 4378
rect 17802 4326 17854 4378
rect 17866 4326 17918 4378
rect 1860 4156 1912 4208
rect 2596 4224 2648 4276
rect 3884 4224 3936 4276
rect 4436 4224 4488 4276
rect 5080 4224 5132 4276
rect 5172 4224 5224 4276
rect 12992 4224 13044 4276
rect 15200 4224 15252 4276
rect 5816 4199 5868 4208
rect 1676 4088 1728 4140
rect 2228 4088 2280 4140
rect 3884 4088 3936 4140
rect 4252 4088 4304 4140
rect 4344 4131 4396 4140
rect 4344 4097 4353 4131
rect 4353 4097 4387 4131
rect 4387 4097 4396 4131
rect 4344 4088 4396 4097
rect 4620 4131 4672 4140
rect 4620 4097 4629 4131
rect 4629 4097 4663 4131
rect 4663 4097 4672 4131
rect 4620 4088 4672 4097
rect 5264 4131 5316 4140
rect 5264 4097 5273 4131
rect 5273 4097 5307 4131
rect 5307 4097 5316 4131
rect 5264 4088 5316 4097
rect 5816 4165 5825 4199
rect 5825 4165 5859 4199
rect 5859 4165 5868 4199
rect 5816 4156 5868 4165
rect 6460 4156 6512 4208
rect 7472 4088 7524 4140
rect 8300 4156 8352 4208
rect 8760 4156 8812 4208
rect 9404 4156 9456 4208
rect 9956 4156 10008 4208
rect 11980 4156 12032 4208
rect 2320 3952 2372 4004
rect 4804 4020 4856 4072
rect 5448 4020 5500 4072
rect 5540 4020 5592 4072
rect 10968 4088 11020 4140
rect 11152 4088 11204 4140
rect 12348 4088 12400 4140
rect 13084 4156 13136 4208
rect 16396 4156 16448 4208
rect 13912 4088 13964 4140
rect 14924 4088 14976 4140
rect 17316 4088 17368 4140
rect 18236 4131 18288 4140
rect 18236 4097 18245 4131
rect 18245 4097 18279 4131
rect 18279 4097 18288 4131
rect 18236 4088 18288 4097
rect 9588 4063 9640 4072
rect 9588 4029 9597 4063
rect 9597 4029 9631 4063
rect 9631 4029 9640 4063
rect 9588 4020 9640 4029
rect 9772 4063 9824 4072
rect 9772 4029 9781 4063
rect 9781 4029 9815 4063
rect 9815 4029 9824 4063
rect 9772 4020 9824 4029
rect 10048 4063 10100 4072
rect 10048 4029 10057 4063
rect 10057 4029 10091 4063
rect 10091 4029 10100 4063
rect 10048 4020 10100 4029
rect 10416 4020 10468 4072
rect 11336 4020 11388 4072
rect 11796 4020 11848 4072
rect 4344 3952 4396 4004
rect 13452 3952 13504 4004
rect 13728 4020 13780 4072
rect 17960 4020 18012 4072
rect 2964 3884 3016 3936
rect 4896 3884 4948 3936
rect 5448 3927 5500 3936
rect 5448 3893 5457 3927
rect 5457 3893 5491 3927
rect 5491 3893 5500 3927
rect 5448 3884 5500 3893
rect 5908 3884 5960 3936
rect 6460 3884 6512 3936
rect 8300 3884 8352 3936
rect 9404 3884 9456 3936
rect 11152 3884 11204 3936
rect 11520 3884 11572 3936
rect 14372 3952 14424 4004
rect 14924 3952 14976 4004
rect 15108 3952 15160 4004
rect 17868 3952 17920 4004
rect 15384 3884 15436 3936
rect 17408 3884 17460 3936
rect 18420 3927 18472 3936
rect 18420 3893 18429 3927
rect 18429 3893 18463 3927
rect 18463 3893 18472 3927
rect 18420 3884 18472 3893
rect 1950 3782 2002 3834
rect 2014 3782 2066 3834
rect 2078 3782 2130 3834
rect 2142 3782 2194 3834
rect 2206 3782 2258 3834
rect 6950 3782 7002 3834
rect 7014 3782 7066 3834
rect 7078 3782 7130 3834
rect 7142 3782 7194 3834
rect 7206 3782 7258 3834
rect 11950 3782 12002 3834
rect 12014 3782 12066 3834
rect 12078 3782 12130 3834
rect 12142 3782 12194 3834
rect 12206 3782 12258 3834
rect 16950 3782 17002 3834
rect 17014 3782 17066 3834
rect 17078 3782 17130 3834
rect 17142 3782 17194 3834
rect 17206 3782 17258 3834
rect 296 3680 348 3732
rect 5448 3680 5500 3732
rect 1032 3612 1084 3664
rect 2320 3612 2372 3664
rect 3056 3612 3108 3664
rect 6368 3680 6420 3732
rect 9680 3680 9732 3732
rect 10232 3680 10284 3732
rect 11428 3680 11480 3732
rect 11704 3680 11756 3732
rect 16396 3680 16448 3732
rect 16580 3680 16632 3732
rect 17868 3723 17920 3732
rect 17868 3689 17877 3723
rect 17877 3689 17911 3723
rect 17911 3689 17920 3723
rect 17868 3680 17920 3689
rect 17960 3680 18012 3732
rect 5632 3612 5684 3664
rect 2872 3544 2924 3596
rect 5816 3544 5868 3596
rect 6552 3544 6604 3596
rect 1400 3519 1452 3528
rect 1400 3485 1409 3519
rect 1409 3485 1443 3519
rect 1443 3485 1452 3519
rect 1400 3476 1452 3485
rect 1860 3476 1912 3528
rect 2688 3519 2740 3528
rect 2688 3485 2697 3519
rect 2697 3485 2731 3519
rect 2731 3485 2740 3519
rect 2688 3476 2740 3485
rect 1400 3340 1452 3392
rect 1952 3340 2004 3392
rect 3056 3519 3108 3528
rect 3056 3485 3065 3519
rect 3065 3485 3099 3519
rect 3099 3485 3108 3519
rect 3056 3476 3108 3485
rect 4160 3519 4212 3528
rect 4160 3485 4169 3519
rect 4169 3485 4203 3519
rect 4203 3485 4212 3519
rect 4160 3476 4212 3485
rect 4344 3519 4396 3528
rect 4344 3485 4353 3519
rect 4353 3485 4387 3519
rect 4387 3485 4396 3519
rect 4344 3476 4396 3485
rect 4528 3519 4580 3528
rect 4528 3485 4537 3519
rect 4537 3485 4571 3519
rect 4571 3485 4580 3519
rect 4528 3476 4580 3485
rect 5264 3476 5316 3528
rect 3240 3408 3292 3460
rect 2964 3340 3016 3392
rect 4896 3408 4948 3460
rect 6092 3476 6144 3528
rect 5540 3408 5592 3460
rect 6920 3476 6972 3528
rect 7012 3519 7064 3528
rect 7288 3544 7340 3596
rect 7012 3485 7061 3519
rect 7061 3485 7064 3519
rect 7012 3476 7064 3485
rect 7380 3476 7432 3528
rect 8116 3544 8168 3596
rect 10876 3612 10928 3664
rect 6368 3451 6420 3460
rect 6368 3417 6377 3451
rect 6377 3417 6411 3451
rect 6411 3417 6420 3451
rect 6368 3408 6420 3417
rect 8208 3519 8260 3528
rect 8208 3485 8217 3519
rect 8217 3485 8251 3519
rect 8251 3485 8260 3519
rect 8208 3476 8260 3485
rect 8300 3519 8352 3528
rect 8300 3485 8309 3519
rect 8309 3485 8343 3519
rect 8343 3485 8352 3519
rect 8300 3476 8352 3485
rect 9680 3544 9732 3596
rect 12808 3612 12860 3664
rect 13176 3612 13228 3664
rect 11796 3544 11848 3596
rect 14004 3544 14056 3596
rect 15292 3544 15344 3596
rect 15752 3544 15804 3596
rect 15936 3587 15988 3596
rect 15936 3553 15945 3587
rect 15945 3553 15979 3587
rect 15979 3553 15988 3587
rect 15936 3544 15988 3553
rect 5632 3340 5684 3392
rect 8484 3408 8536 3460
rect 8760 3451 8812 3460
rect 8760 3417 8769 3451
rect 8769 3417 8803 3451
rect 8803 3417 8812 3451
rect 8760 3408 8812 3417
rect 9220 3476 9272 3528
rect 9312 3519 9364 3528
rect 9312 3485 9321 3519
rect 9321 3485 9355 3519
rect 9355 3485 9364 3519
rect 9312 3476 9364 3485
rect 9496 3476 9548 3528
rect 11888 3476 11940 3528
rect 12624 3519 12676 3528
rect 12624 3485 12633 3519
rect 12633 3485 12667 3519
rect 12667 3485 12676 3519
rect 12624 3476 12676 3485
rect 12716 3519 12768 3528
rect 12716 3485 12725 3519
rect 12725 3485 12759 3519
rect 12759 3485 12768 3519
rect 12716 3476 12768 3485
rect 13452 3476 13504 3528
rect 13636 3476 13688 3528
rect 9864 3408 9916 3460
rect 8024 3340 8076 3392
rect 8208 3340 8260 3392
rect 8852 3340 8904 3392
rect 10876 3408 10928 3460
rect 12072 3340 12124 3392
rect 12532 3340 12584 3392
rect 12624 3340 12676 3392
rect 13360 3340 13412 3392
rect 15384 3451 15436 3460
rect 15384 3417 15393 3451
rect 15393 3417 15427 3451
rect 15427 3417 15436 3451
rect 15384 3408 15436 3417
rect 16028 3519 16080 3528
rect 16028 3485 16037 3519
rect 16037 3485 16071 3519
rect 16071 3485 16080 3519
rect 16028 3476 16080 3485
rect 16396 3519 16448 3528
rect 16396 3485 16405 3519
rect 16405 3485 16439 3519
rect 16439 3485 16448 3519
rect 16396 3476 16448 3485
rect 16304 3408 16356 3460
rect 16580 3476 16632 3528
rect 16856 3519 16908 3528
rect 16856 3485 16865 3519
rect 16865 3485 16899 3519
rect 16899 3485 16908 3519
rect 16856 3476 16908 3485
rect 17408 3587 17460 3596
rect 17408 3553 17417 3587
rect 17417 3553 17451 3587
rect 17451 3553 17460 3587
rect 17408 3544 17460 3553
rect 17316 3519 17368 3528
rect 17316 3485 17325 3519
rect 17325 3485 17359 3519
rect 17359 3485 17368 3519
rect 17316 3476 17368 3485
rect 17500 3476 17552 3528
rect 18052 3544 18104 3596
rect 17960 3519 18012 3528
rect 17960 3485 17969 3519
rect 17969 3485 18003 3519
rect 18003 3485 18012 3519
rect 17960 3476 18012 3485
rect 18144 3519 18196 3528
rect 18144 3485 18153 3519
rect 18153 3485 18187 3519
rect 18187 3485 18196 3519
rect 18144 3476 18196 3485
rect 2610 3238 2662 3290
rect 2674 3238 2726 3290
rect 2738 3238 2790 3290
rect 2802 3238 2854 3290
rect 2866 3238 2918 3290
rect 7610 3238 7662 3290
rect 7674 3238 7726 3290
rect 7738 3238 7790 3290
rect 7802 3238 7854 3290
rect 7866 3238 7918 3290
rect 12610 3238 12662 3290
rect 12674 3238 12726 3290
rect 12738 3238 12790 3290
rect 12802 3238 12854 3290
rect 12866 3238 12918 3290
rect 17610 3238 17662 3290
rect 17674 3238 17726 3290
rect 17738 3238 17790 3290
rect 17802 3238 17854 3290
rect 17866 3238 17918 3290
rect 3700 3136 3752 3188
rect 6736 3136 6788 3188
rect 7472 3136 7524 3188
rect 8944 3179 8996 3188
rect 8944 3145 8953 3179
rect 8953 3145 8987 3179
rect 8987 3145 8996 3179
rect 8944 3136 8996 3145
rect 5172 3068 5224 3120
rect 5448 3068 5500 3120
rect 2412 3043 2464 3052
rect 2412 3009 2421 3043
rect 2421 3009 2455 3043
rect 2455 3009 2464 3043
rect 2412 3000 2464 3009
rect 2780 3043 2832 3052
rect 2780 3009 2789 3043
rect 2789 3009 2823 3043
rect 2823 3009 2832 3043
rect 2780 3000 2832 3009
rect 2964 3043 3016 3052
rect 2964 3009 2973 3043
rect 2973 3009 3007 3043
rect 3007 3009 3016 3043
rect 2964 3000 3016 3009
rect 3332 3000 3384 3052
rect 3516 3043 3568 3052
rect 3516 3009 3525 3043
rect 3525 3009 3559 3043
rect 3559 3009 3568 3043
rect 3516 3000 3568 3009
rect 2504 2932 2556 2984
rect 3148 2975 3200 2984
rect 3148 2941 3157 2975
rect 3157 2941 3191 2975
rect 3191 2941 3200 2975
rect 3148 2932 3200 2941
rect 3240 2975 3292 2984
rect 3240 2941 3249 2975
rect 3249 2941 3283 2975
rect 3283 2941 3292 2975
rect 3240 2932 3292 2941
rect 5724 3000 5776 3052
rect 4252 2932 4304 2984
rect 7656 3068 7708 3120
rect 6552 3043 6604 3052
rect 6552 3009 6561 3043
rect 6561 3009 6595 3043
rect 6595 3009 6604 3043
rect 6552 3000 6604 3009
rect 6644 3000 6696 3052
rect 6460 2932 6512 2984
rect 8300 3043 8352 3052
rect 8300 3009 8309 3043
rect 8309 3009 8343 3043
rect 8343 3009 8352 3043
rect 8300 3000 8352 3009
rect 8392 3065 8444 3074
rect 8392 3031 8401 3065
rect 8401 3031 8435 3065
rect 8435 3031 8444 3065
rect 8392 3022 8444 3031
rect 9128 3068 9180 3120
rect 3884 2907 3936 2916
rect 3884 2873 3893 2907
rect 3893 2873 3927 2907
rect 3927 2873 3936 2907
rect 3884 2864 3936 2873
rect 5080 2864 5132 2916
rect 7932 2975 7984 2984
rect 7932 2941 7941 2975
rect 7941 2941 7975 2975
rect 7975 2941 7984 2975
rect 7932 2932 7984 2941
rect 8576 2975 8628 2984
rect 8576 2941 8585 2975
rect 8585 2941 8619 2975
rect 8619 2941 8628 2975
rect 8576 2932 8628 2941
rect 8852 2932 8904 2984
rect 9312 3043 9364 3052
rect 9312 3009 9321 3043
rect 9321 3009 9355 3043
rect 9355 3009 9364 3043
rect 9312 3000 9364 3009
rect 10416 3136 10468 3188
rect 11704 3179 11756 3188
rect 11704 3145 11731 3179
rect 11731 3145 11756 3179
rect 11704 3136 11756 3145
rect 14096 3136 14148 3188
rect 14464 3136 14516 3188
rect 17408 3136 17460 3188
rect 9956 3068 10008 3120
rect 11060 3068 11112 3120
rect 11888 3111 11940 3120
rect 11888 3077 11897 3111
rect 11897 3077 11931 3111
rect 11931 3077 11940 3111
rect 11888 3068 11940 3077
rect 9588 3043 9640 3052
rect 9588 3009 9597 3043
rect 9597 3009 9631 3043
rect 9631 3009 9640 3043
rect 9588 3000 9640 3009
rect 10784 3000 10836 3052
rect 10968 3000 11020 3052
rect 11612 3000 11664 3052
rect 16212 3068 16264 3120
rect 12072 3043 12124 3052
rect 12072 3009 12081 3043
rect 12081 3009 12115 3043
rect 12115 3009 12124 3043
rect 12072 3000 12124 3009
rect 11244 2932 11296 2984
rect 12440 3000 12492 3052
rect 12716 2975 12768 2984
rect 12716 2941 12725 2975
rect 12725 2941 12759 2975
rect 12759 2941 12768 2975
rect 12716 2932 12768 2941
rect 13084 3043 13136 3052
rect 13084 3009 13093 3043
rect 13093 3009 13127 3043
rect 13127 3009 13136 3043
rect 13084 3000 13136 3009
rect 13636 3000 13688 3052
rect 15844 3000 15896 3052
rect 16488 3000 16540 3052
rect 16948 2932 17000 2984
rect 17316 2932 17368 2984
rect 6644 2907 6696 2916
rect 6644 2873 6653 2907
rect 6653 2873 6687 2907
rect 6687 2873 6696 2907
rect 6644 2864 6696 2873
rect 6736 2907 6788 2916
rect 6736 2873 6745 2907
rect 6745 2873 6779 2907
rect 6779 2873 6788 2907
rect 6736 2864 6788 2873
rect 2964 2796 3016 2848
rect 3976 2839 4028 2848
rect 3976 2805 3985 2839
rect 3985 2805 4019 2839
rect 4019 2805 4028 2839
rect 3976 2796 4028 2805
rect 4896 2796 4948 2848
rect 6552 2796 6604 2848
rect 7840 2796 7892 2848
rect 8208 2864 8260 2916
rect 10600 2796 10652 2848
rect 10784 2796 10836 2848
rect 11336 2796 11388 2848
rect 11612 2796 11664 2848
rect 12348 2864 12400 2916
rect 13360 2864 13412 2916
rect 18052 2864 18104 2916
rect 14188 2796 14240 2848
rect 16856 2796 16908 2848
rect 1950 2694 2002 2746
rect 2014 2694 2066 2746
rect 2078 2694 2130 2746
rect 2142 2694 2194 2746
rect 2206 2694 2258 2746
rect 6950 2694 7002 2746
rect 7014 2694 7066 2746
rect 7078 2694 7130 2746
rect 7142 2694 7194 2746
rect 7206 2694 7258 2746
rect 11950 2694 12002 2746
rect 12014 2694 12066 2746
rect 12078 2694 12130 2746
rect 12142 2694 12194 2746
rect 12206 2694 12258 2746
rect 16950 2694 17002 2746
rect 17014 2694 17066 2746
rect 17078 2694 17130 2746
rect 17142 2694 17194 2746
rect 17206 2694 17258 2746
rect 1676 2592 1728 2644
rect 3424 2592 3476 2644
rect 3792 2592 3844 2644
rect 5448 2592 5500 2644
rect 9036 2635 9088 2644
rect 9036 2601 9045 2635
rect 9045 2601 9079 2635
rect 9079 2601 9088 2635
rect 9036 2592 9088 2601
rect 9220 2592 9272 2644
rect 480 2456 532 2508
rect 1308 2388 1360 2440
rect 1676 2388 1728 2440
rect 1860 2431 1912 2440
rect 1860 2397 1869 2431
rect 1869 2397 1903 2431
rect 1903 2397 1912 2431
rect 1860 2388 1912 2397
rect 4988 2456 5040 2508
rect 6552 2524 6604 2576
rect 9312 2524 9364 2576
rect 13360 2592 13412 2644
rect 11428 2524 11480 2576
rect 6736 2456 6788 2508
rect 7472 2456 7524 2508
rect 2044 2431 2096 2440
rect 2044 2397 2053 2431
rect 2053 2397 2087 2431
rect 2087 2397 2096 2431
rect 2044 2388 2096 2397
rect 2412 2388 2464 2440
rect 4252 2388 4304 2440
rect 6552 2431 6604 2440
rect 6552 2397 6561 2431
rect 6561 2397 6595 2431
rect 6595 2397 6604 2431
rect 6552 2388 6604 2397
rect 8484 2456 8536 2508
rect 8576 2499 8628 2508
rect 8576 2465 8585 2499
rect 8585 2465 8619 2499
rect 8619 2465 8628 2499
rect 8576 2456 8628 2465
rect 8668 2499 8720 2508
rect 8668 2465 8677 2499
rect 8677 2465 8711 2499
rect 8711 2465 8720 2499
rect 8668 2456 8720 2465
rect 9404 2456 9456 2508
rect 11060 2456 11112 2508
rect 13820 2456 13872 2508
rect 15292 2456 15344 2508
rect 18512 2456 18564 2508
rect 8760 2388 8812 2440
rect 9220 2431 9272 2440
rect 9220 2397 9229 2431
rect 9229 2397 9263 2431
rect 9263 2397 9272 2431
rect 9220 2388 9272 2397
rect 9312 2431 9364 2440
rect 9312 2397 9321 2431
rect 9321 2397 9355 2431
rect 9355 2397 9364 2431
rect 9312 2388 9364 2397
rect 9588 2431 9640 2440
rect 9588 2397 9597 2431
rect 9597 2397 9631 2431
rect 9631 2397 9640 2431
rect 9588 2388 9640 2397
rect 3332 2320 3384 2372
rect 8208 2320 8260 2372
rect 10876 2388 10928 2440
rect 11152 2431 11204 2440
rect 11152 2397 11161 2431
rect 11161 2397 11195 2431
rect 11195 2397 11204 2431
rect 11152 2388 11204 2397
rect 11336 2431 11388 2440
rect 11336 2397 11345 2431
rect 11345 2397 11379 2431
rect 11379 2397 11388 2431
rect 11336 2388 11388 2397
rect 11612 2388 11664 2440
rect 11704 2388 11756 2440
rect 11980 2431 12032 2440
rect 11980 2397 11989 2431
rect 11989 2397 12023 2431
rect 12023 2397 12032 2431
rect 11980 2388 12032 2397
rect 12440 2388 12492 2440
rect 12808 2388 12860 2440
rect 13728 2388 13780 2440
rect 16580 2388 16632 2440
rect 16948 2388 17000 2440
rect 9956 2320 10008 2372
rect 15660 2320 15712 2372
rect 18328 2363 18380 2372
rect 18328 2329 18337 2363
rect 18337 2329 18371 2363
rect 18371 2329 18380 2363
rect 18328 2320 18380 2329
rect 2504 2295 2556 2304
rect 2504 2261 2513 2295
rect 2513 2261 2547 2295
rect 2547 2261 2556 2295
rect 2504 2252 2556 2261
rect 4528 2252 4580 2304
rect 7196 2295 7248 2304
rect 7196 2261 7205 2295
rect 7205 2261 7239 2295
rect 7239 2261 7248 2295
rect 7196 2252 7248 2261
rect 7656 2252 7708 2304
rect 9128 2252 9180 2304
rect 11060 2252 11112 2304
rect 11612 2295 11664 2304
rect 11612 2261 11621 2295
rect 11621 2261 11655 2295
rect 11655 2261 11664 2295
rect 11612 2252 11664 2261
rect 12440 2252 12492 2304
rect 13268 2252 13320 2304
rect 16856 2295 16908 2304
rect 16856 2261 16865 2295
rect 16865 2261 16899 2295
rect 16899 2261 16908 2295
rect 16856 2252 16908 2261
rect 2610 2150 2662 2202
rect 2674 2150 2726 2202
rect 2738 2150 2790 2202
rect 2802 2150 2854 2202
rect 2866 2150 2918 2202
rect 7610 2150 7662 2202
rect 7674 2150 7726 2202
rect 7738 2150 7790 2202
rect 7802 2150 7854 2202
rect 7866 2150 7918 2202
rect 12610 2150 12662 2202
rect 12674 2150 12726 2202
rect 12738 2150 12790 2202
rect 12802 2150 12854 2202
rect 12866 2150 12918 2202
rect 17610 2150 17662 2202
rect 17674 2150 17726 2202
rect 17738 2150 17790 2202
rect 17802 2150 17854 2202
rect 17866 2150 17918 2202
rect 6736 2048 6788 2100
rect 9404 2048 9456 2100
rect 10784 2048 10836 2100
rect 13176 2048 13228 2100
rect 848 1980 900 2032
rect 9220 1980 9272 2032
rect 10968 1980 11020 2032
rect 13544 1980 13596 2032
rect 16856 1980 16908 2032
rect 4068 1912 4120 1964
rect 10692 1912 10744 1964
rect 9312 1844 9364 1896
rect 17960 1844 18012 1896
rect 3056 1776 3108 1828
rect 11520 1776 11572 1828
rect 7472 1708 7524 1760
rect 11060 1708 11112 1760
rect 1676 1640 1728 1692
rect 6460 1640 6512 1692
rect 14924 1708 14976 1760
rect 6276 1572 6328 1624
rect 9772 1572 9824 1624
rect 8484 1504 8536 1556
rect 17500 1504 17552 1556
rect 5724 1436 5776 1488
rect 13084 1436 13136 1488
rect 2320 1300 2372 1352
rect 6092 1300 6144 1352
rect 6184 1300 6236 1352
rect 11152 1300 11204 1352
rect 4620 1232 4672 1284
rect 11244 1232 11296 1284
rect 7288 1164 7340 1216
rect 12992 1232 13044 1284
rect 6368 1096 6420 1148
rect 16764 1164 16816 1216
rect 2964 1028 3016 1080
rect 5816 1028 5868 1080
rect 16028 1028 16080 1080
rect 4160 960 4212 1012
rect 11796 960 11848 1012
rect 3148 892 3200 944
rect 15384 892 15436 944
rect 6000 824 6052 876
rect 15476 824 15528 876
rect 5172 756 5224 808
rect 17316 756 17368 808
rect 5264 620 5316 672
rect 12532 620 12584 672
rect 6644 552 6696 604
rect 14280 552 14332 604
rect 3976 484 4028 536
rect 14648 484 14700 536
<< metal2 >>
rect 1214 19200 1270 20000
rect 3698 19200 3754 20000
rect 6182 19200 6238 20000
rect 8666 19200 8722 20000
rect 11150 19200 11206 20000
rect 13634 19200 13690 20000
rect 16118 19200 16174 20000
rect 18602 19200 18658 20000
rect 1122 18728 1178 18737
rect 1122 18663 1178 18672
rect 754 17776 810 17785
rect 754 17711 810 17720
rect 204 15496 256 15502
rect 204 15438 256 15444
rect 110 12336 166 12345
rect 110 12271 166 12280
rect 124 9722 152 12271
rect 112 9716 164 9722
rect 112 9658 164 9664
rect 124 7002 152 9658
rect 216 8430 244 15438
rect 296 13796 348 13802
rect 296 13738 348 13744
rect 204 8424 256 8430
rect 204 8366 256 8372
rect 112 6996 164 7002
rect 112 6938 164 6944
rect 308 3738 336 13738
rect 480 12776 532 12782
rect 480 12718 532 12724
rect 388 9580 440 9586
rect 388 9522 440 9528
rect 400 6905 428 9522
rect 386 6896 442 6905
rect 386 6831 442 6840
rect 296 3732 348 3738
rect 296 3674 348 3680
rect 492 2514 520 12718
rect 572 11552 624 11558
rect 572 11494 624 11500
rect 584 6186 612 11494
rect 768 10169 796 17711
rect 940 17332 992 17338
rect 940 17274 992 17280
rect 952 16574 980 17274
rect 952 16546 1072 16574
rect 848 15972 900 15978
rect 848 15914 900 15920
rect 754 10160 810 10169
rect 754 10095 810 10104
rect 754 9072 810 9081
rect 754 9007 810 9016
rect 768 8906 796 9007
rect 756 8900 808 8906
rect 756 8842 808 8848
rect 756 8016 808 8022
rect 756 7958 808 7964
rect 572 6180 624 6186
rect 572 6122 624 6128
rect 768 5642 796 7958
rect 860 7313 888 15914
rect 940 13388 992 13394
rect 940 13330 992 13336
rect 846 7304 902 7313
rect 846 7239 902 7248
rect 848 5772 900 5778
rect 848 5714 900 5720
rect 756 5636 808 5642
rect 756 5578 808 5584
rect 480 2508 532 2514
rect 480 2450 532 2456
rect 860 2038 888 5714
rect 952 3641 980 13330
rect 1044 12457 1072 16546
rect 1136 15094 1164 18663
rect 1228 16590 1256 19200
rect 1584 18624 1636 18630
rect 1584 18566 1636 18572
rect 2962 18592 3018 18601
rect 1306 18320 1362 18329
rect 1306 18255 1362 18264
rect 1216 16584 1268 16590
rect 1216 16526 1268 16532
rect 1320 15162 1348 18255
rect 1492 16516 1544 16522
rect 1492 16458 1544 16464
rect 1504 16153 1532 16458
rect 1490 16144 1546 16153
rect 1490 16079 1546 16088
rect 1400 15428 1452 15434
rect 1400 15370 1452 15376
rect 1308 15156 1360 15162
rect 1308 15098 1360 15104
rect 1124 15088 1176 15094
rect 1124 15030 1176 15036
rect 1412 12458 1440 15370
rect 1596 15337 1624 18566
rect 2962 18527 3018 18536
rect 2318 17640 2374 17649
rect 2318 17575 2374 17584
rect 1768 16992 1820 16998
rect 1768 16934 1820 16940
rect 1780 16017 1808 16934
rect 1950 16892 2258 16901
rect 1950 16890 1956 16892
rect 2012 16890 2036 16892
rect 2092 16890 2116 16892
rect 2172 16890 2196 16892
rect 2252 16890 2258 16892
rect 2012 16838 2014 16890
rect 2194 16838 2196 16890
rect 1950 16836 1956 16838
rect 2012 16836 2036 16838
rect 2092 16836 2116 16838
rect 2172 16836 2196 16838
rect 2252 16836 2258 16838
rect 1950 16827 2258 16836
rect 1860 16652 1912 16658
rect 1860 16594 1912 16600
rect 1766 16008 1822 16017
rect 1766 15943 1822 15952
rect 1872 15858 1900 16594
rect 1780 15830 1900 15858
rect 1582 15328 1638 15337
rect 1582 15263 1638 15272
rect 1780 15178 1808 15830
rect 1950 15804 2258 15813
rect 1950 15802 1956 15804
rect 2012 15802 2036 15804
rect 2092 15802 2116 15804
rect 2172 15802 2196 15804
rect 2252 15802 2258 15804
rect 2012 15750 2014 15802
rect 2194 15750 2196 15802
rect 1950 15748 1956 15750
rect 2012 15748 2036 15750
rect 2092 15748 2116 15750
rect 2172 15748 2196 15750
rect 2252 15748 2258 15750
rect 1950 15739 2258 15748
rect 1860 15700 1912 15706
rect 1860 15642 1912 15648
rect 1596 15150 1808 15178
rect 1492 13932 1544 13938
rect 1492 13874 1544 13880
rect 1504 13705 1532 13874
rect 1490 13696 1546 13705
rect 1490 13631 1546 13640
rect 1596 13546 1624 15150
rect 1768 14952 1820 14958
rect 1768 14894 1820 14900
rect 1780 14618 1808 14894
rect 1768 14612 1820 14618
rect 1768 14554 1820 14560
rect 1872 14482 1900 15642
rect 2332 14958 2360 17575
rect 2610 17436 2918 17445
rect 2610 17434 2616 17436
rect 2672 17434 2696 17436
rect 2752 17434 2776 17436
rect 2832 17434 2856 17436
rect 2912 17434 2918 17436
rect 2672 17382 2674 17434
rect 2854 17382 2856 17434
rect 2610 17380 2616 17382
rect 2672 17380 2696 17382
rect 2752 17380 2776 17382
rect 2832 17380 2856 17382
rect 2912 17380 2918 17382
rect 2610 17371 2918 17380
rect 2976 17270 3004 18527
rect 3332 18488 3384 18494
rect 3332 18430 3384 18436
rect 2964 17264 3016 17270
rect 2964 17206 3016 17212
rect 3056 17196 3108 17202
rect 3056 17138 3108 17144
rect 2412 16992 2464 16998
rect 2410 16960 2412 16969
rect 2464 16960 2466 16969
rect 2410 16895 2466 16904
rect 2610 16348 2918 16357
rect 2610 16346 2616 16348
rect 2672 16346 2696 16348
rect 2752 16346 2776 16348
rect 2832 16346 2856 16348
rect 2912 16346 2918 16348
rect 2672 16294 2674 16346
rect 2854 16294 2856 16346
rect 2610 16292 2616 16294
rect 2672 16292 2696 16294
rect 2752 16292 2776 16294
rect 2832 16292 2856 16294
rect 2912 16292 2918 16294
rect 2610 16283 2918 16292
rect 3068 16114 3096 17138
rect 3148 16516 3200 16522
rect 3148 16458 3200 16464
rect 3056 16108 3108 16114
rect 2976 16068 3056 16096
rect 2780 16040 2832 16046
rect 2780 15982 2832 15988
rect 2792 15638 2820 15982
rect 2780 15632 2832 15638
rect 2502 15600 2558 15609
rect 2780 15574 2832 15580
rect 2502 15535 2558 15544
rect 2412 15360 2464 15366
rect 2412 15302 2464 15308
rect 2320 14952 2372 14958
rect 2320 14894 2372 14900
rect 1950 14716 2258 14725
rect 1950 14714 1956 14716
rect 2012 14714 2036 14716
rect 2092 14714 2116 14716
rect 2172 14714 2196 14716
rect 2252 14714 2258 14716
rect 2012 14662 2014 14714
rect 2194 14662 2196 14714
rect 1950 14660 1956 14662
rect 2012 14660 2036 14662
rect 2092 14660 2116 14662
rect 2172 14660 2196 14662
rect 2252 14660 2258 14662
rect 1950 14651 2258 14660
rect 2228 14612 2280 14618
rect 2228 14554 2280 14560
rect 2240 14482 2268 14554
rect 1676 14476 1728 14482
rect 1676 14418 1728 14424
rect 1860 14476 1912 14482
rect 1860 14418 1912 14424
rect 2228 14476 2280 14482
rect 2228 14418 2280 14424
rect 1030 12448 1086 12457
rect 1320 12434 1440 12458
rect 1030 12383 1086 12392
rect 1228 12430 1440 12434
rect 1504 13518 1624 13546
rect 1228 12406 1348 12430
rect 1228 12288 1256 12406
rect 1044 12260 1256 12288
rect 1308 12300 1360 12306
rect 1044 9761 1072 12260
rect 1308 12242 1360 12248
rect 1214 12200 1270 12209
rect 1214 12135 1270 12144
rect 1122 10976 1178 10985
rect 1122 10911 1178 10920
rect 1030 9752 1086 9761
rect 1030 9687 1086 9696
rect 1032 9648 1084 9654
rect 1032 9590 1084 9596
rect 1044 3670 1072 9590
rect 1136 8838 1164 10911
rect 1228 10062 1256 12135
rect 1216 10056 1268 10062
rect 1216 9998 1268 10004
rect 1216 9920 1268 9926
rect 1216 9862 1268 9868
rect 1124 8832 1176 8838
rect 1124 8774 1176 8780
rect 1124 8628 1176 8634
rect 1124 8570 1176 8576
rect 1136 5370 1164 8570
rect 1124 5364 1176 5370
rect 1124 5306 1176 5312
rect 1228 4049 1256 9862
rect 1320 8401 1348 12242
rect 1400 12232 1452 12238
rect 1400 12174 1452 12180
rect 1412 11354 1440 12174
rect 1504 11665 1532 13518
rect 1490 11656 1546 11665
rect 1490 11591 1546 11600
rect 1504 11558 1532 11591
rect 1492 11552 1544 11558
rect 1492 11494 1544 11500
rect 1400 11348 1452 11354
rect 1400 11290 1452 11296
rect 1584 11280 1636 11286
rect 1398 11248 1454 11257
rect 1584 11222 1636 11228
rect 1398 11183 1454 11192
rect 1492 11212 1544 11218
rect 1412 11150 1440 11183
rect 1492 11154 1544 11160
rect 1400 11144 1452 11150
rect 1400 11086 1452 11092
rect 1400 11008 1452 11014
rect 1400 10950 1452 10956
rect 1412 10266 1440 10950
rect 1400 10260 1452 10266
rect 1400 10202 1452 10208
rect 1400 10056 1452 10062
rect 1400 9998 1452 10004
rect 1306 8392 1362 8401
rect 1306 8327 1362 8336
rect 1308 7744 1360 7750
rect 1308 7686 1360 7692
rect 1320 5574 1348 7686
rect 1412 5846 1440 9998
rect 1504 7478 1532 11154
rect 1596 9654 1624 11222
rect 1688 10130 1716 14418
rect 1952 14408 2004 14414
rect 1858 14376 1914 14385
rect 1952 14350 2004 14356
rect 2136 14408 2188 14414
rect 2136 14350 2188 14356
rect 1858 14311 1914 14320
rect 1768 13184 1820 13190
rect 1768 13126 1820 13132
rect 1780 11218 1808 13126
rect 1872 12782 1900 14311
rect 1964 13977 1992 14350
rect 2148 14249 2176 14350
rect 2134 14240 2190 14249
rect 2134 14175 2190 14184
rect 1950 13968 2006 13977
rect 1950 13903 2006 13912
rect 1950 13628 2258 13637
rect 1950 13626 1956 13628
rect 2012 13626 2036 13628
rect 2092 13626 2116 13628
rect 2172 13626 2196 13628
rect 2252 13626 2258 13628
rect 2012 13574 2014 13626
rect 2194 13574 2196 13626
rect 1950 13572 1956 13574
rect 2012 13572 2036 13574
rect 2092 13572 2116 13574
rect 2172 13572 2196 13574
rect 2252 13572 2258 13574
rect 1950 13563 2258 13572
rect 2228 13524 2280 13530
rect 2228 13466 2280 13472
rect 2240 12918 2268 13466
rect 2320 13320 2372 13326
rect 2320 13262 2372 13268
rect 2332 12986 2360 13262
rect 2320 12980 2372 12986
rect 2320 12922 2372 12928
rect 1952 12912 2004 12918
rect 1952 12854 2004 12860
rect 2228 12912 2280 12918
rect 2228 12854 2280 12860
rect 1860 12776 1912 12782
rect 1860 12718 1912 12724
rect 1964 12628 1992 12854
rect 1872 12600 1992 12628
rect 1872 11558 1900 12600
rect 1950 12540 2258 12549
rect 1950 12538 1956 12540
rect 2012 12538 2036 12540
rect 2092 12538 2116 12540
rect 2172 12538 2196 12540
rect 2252 12538 2258 12540
rect 2012 12486 2014 12538
rect 2194 12486 2196 12538
rect 1950 12484 1956 12486
rect 2012 12484 2036 12486
rect 2092 12484 2116 12486
rect 2172 12484 2196 12486
rect 2252 12484 2258 12486
rect 1950 12475 2258 12484
rect 2136 12436 2188 12442
rect 2424 12424 2452 15302
rect 2516 13814 2544 15535
rect 2610 15260 2918 15269
rect 2610 15258 2616 15260
rect 2672 15258 2696 15260
rect 2752 15258 2776 15260
rect 2832 15258 2856 15260
rect 2912 15258 2918 15260
rect 2672 15206 2674 15258
rect 2854 15206 2856 15258
rect 2610 15204 2616 15206
rect 2672 15204 2696 15206
rect 2752 15204 2776 15206
rect 2832 15204 2856 15206
rect 2912 15204 2918 15206
rect 2610 15195 2918 15204
rect 2976 14482 3004 16068
rect 3056 16050 3108 16056
rect 3160 15008 3188 16458
rect 3240 15632 3292 15638
rect 3240 15574 3292 15580
rect 3068 14980 3188 15008
rect 2964 14476 3016 14482
rect 2964 14418 3016 14424
rect 2610 14172 2918 14181
rect 2610 14170 2616 14172
rect 2672 14170 2696 14172
rect 2752 14170 2776 14172
rect 2832 14170 2856 14172
rect 2912 14170 2918 14172
rect 2672 14118 2674 14170
rect 2854 14118 2856 14170
rect 2610 14116 2616 14118
rect 2672 14116 2696 14118
rect 2752 14116 2776 14118
rect 2832 14116 2856 14118
rect 2912 14116 2918 14118
rect 2610 14107 2918 14116
rect 2872 14068 2924 14074
rect 2872 14010 2924 14016
rect 2884 13938 2912 14010
rect 2976 13938 3004 14418
rect 2872 13932 2924 13938
rect 2872 13874 2924 13880
rect 2964 13932 3016 13938
rect 2964 13874 3016 13880
rect 2516 13786 2636 13814
rect 2608 13326 2636 13786
rect 2504 13320 2556 13326
rect 2504 13262 2556 13268
rect 2596 13320 2648 13326
rect 2872 13320 2924 13326
rect 2596 13262 2648 13268
rect 2870 13288 2872 13297
rect 2964 13320 3016 13326
rect 2924 13288 2926 13297
rect 2516 12866 2544 13262
rect 2964 13262 3016 13268
rect 2870 13223 2926 13232
rect 2610 13084 2918 13093
rect 2610 13082 2616 13084
rect 2672 13082 2696 13084
rect 2752 13082 2776 13084
rect 2832 13082 2856 13084
rect 2912 13082 2918 13084
rect 2672 13030 2674 13082
rect 2854 13030 2856 13082
rect 2610 13028 2616 13030
rect 2672 13028 2696 13030
rect 2752 13028 2776 13030
rect 2832 13028 2856 13030
rect 2912 13028 2918 13030
rect 2610 13019 2918 13028
rect 2976 12986 3004 13262
rect 2688 12980 2740 12986
rect 2688 12922 2740 12928
rect 2964 12980 3016 12986
rect 2964 12922 3016 12928
rect 2516 12838 2636 12866
rect 2504 12776 2556 12782
rect 2504 12718 2556 12724
rect 2136 12378 2188 12384
rect 2332 12396 2452 12424
rect 2148 11558 2176 12378
rect 1860 11552 1912 11558
rect 1860 11494 1912 11500
rect 2136 11552 2188 11558
rect 2136 11494 2188 11500
rect 1768 11212 1820 11218
rect 1768 11154 1820 11160
rect 1768 11076 1820 11082
rect 1768 11018 1820 11024
rect 1676 10124 1728 10130
rect 1676 10066 1728 10072
rect 1584 9648 1636 9654
rect 1584 9590 1636 9596
rect 1676 9376 1728 9382
rect 1676 9318 1728 9324
rect 1582 9072 1638 9081
rect 1582 9007 1638 9016
rect 1596 8974 1624 9007
rect 1584 8968 1636 8974
rect 1584 8910 1636 8916
rect 1584 8832 1636 8838
rect 1584 8774 1636 8780
rect 1492 7472 1544 7478
rect 1492 7414 1544 7420
rect 1492 6724 1544 6730
rect 1492 6666 1544 6672
rect 1504 6361 1532 6666
rect 1490 6352 1546 6361
rect 1490 6287 1546 6296
rect 1596 6236 1624 8774
rect 1688 8634 1716 9318
rect 1676 8628 1728 8634
rect 1676 8570 1728 8576
rect 1780 8566 1808 11018
rect 1872 10198 1900 11494
rect 1950 11452 2258 11461
rect 1950 11450 1956 11452
rect 2012 11450 2036 11452
rect 2092 11450 2116 11452
rect 2172 11450 2196 11452
rect 2252 11450 2258 11452
rect 2012 11398 2014 11450
rect 2194 11398 2196 11450
rect 1950 11396 1956 11398
rect 2012 11396 2036 11398
rect 2092 11396 2116 11398
rect 2172 11396 2196 11398
rect 2252 11396 2258 11398
rect 1950 11387 2258 11396
rect 2228 11348 2280 11354
rect 2228 11290 2280 11296
rect 2240 10810 2268 11290
rect 2228 10804 2280 10810
rect 2228 10746 2280 10752
rect 1950 10364 2258 10373
rect 1950 10362 1956 10364
rect 2012 10362 2036 10364
rect 2092 10362 2116 10364
rect 2172 10362 2196 10364
rect 2252 10362 2258 10364
rect 2012 10310 2014 10362
rect 2194 10310 2196 10362
rect 1950 10308 1956 10310
rect 2012 10308 2036 10310
rect 2092 10308 2116 10310
rect 2172 10308 2196 10310
rect 2252 10308 2258 10310
rect 1950 10299 2258 10308
rect 1952 10260 2004 10266
rect 1952 10202 2004 10208
rect 1860 10192 1912 10198
rect 1860 10134 1912 10140
rect 1964 9466 1992 10202
rect 2136 10192 2188 10198
rect 2136 10134 2188 10140
rect 2228 10192 2280 10198
rect 2228 10134 2280 10140
rect 2044 9580 2096 9586
rect 2044 9522 2096 9528
rect 2056 9489 2084 9522
rect 1872 9438 1992 9466
rect 2042 9480 2098 9489
rect 1872 9058 1900 9438
rect 2148 9450 2176 10134
rect 2042 9415 2098 9424
rect 2136 9444 2188 9450
rect 2136 9386 2188 9392
rect 2240 9382 2268 10134
rect 2228 9376 2280 9382
rect 2228 9318 2280 9324
rect 1950 9276 2258 9285
rect 1950 9274 1956 9276
rect 2012 9274 2036 9276
rect 2092 9274 2116 9276
rect 2172 9274 2196 9276
rect 2252 9274 2258 9276
rect 2012 9222 2014 9274
rect 2194 9222 2196 9274
rect 1950 9220 1956 9222
rect 2012 9220 2036 9222
rect 2092 9220 2116 9222
rect 2172 9220 2196 9222
rect 2252 9220 2258 9222
rect 1950 9211 2258 9220
rect 1872 9030 2084 9058
rect 1952 8968 2004 8974
rect 1952 8910 2004 8916
rect 1860 8832 1912 8838
rect 1964 8809 1992 8910
rect 1860 8774 1912 8780
rect 1950 8800 2006 8809
rect 1768 8560 1820 8566
rect 1768 8502 1820 8508
rect 1676 8492 1728 8498
rect 1676 8434 1728 8440
rect 1504 6208 1624 6236
rect 1400 5840 1452 5846
rect 1400 5782 1452 5788
rect 1504 5658 1532 6208
rect 1584 6112 1636 6118
rect 1584 6054 1636 6060
rect 1412 5630 1532 5658
rect 1308 5568 1360 5574
rect 1308 5510 1360 5516
rect 1308 5364 1360 5370
rect 1308 5306 1360 5312
rect 1214 4040 1270 4049
rect 1214 3975 1270 3984
rect 1032 3664 1084 3670
rect 938 3632 994 3641
rect 1032 3606 1084 3612
rect 938 3567 994 3576
rect 1320 2446 1348 5306
rect 1412 4185 1440 5630
rect 1492 5568 1544 5574
rect 1492 5510 1544 5516
rect 1398 4176 1454 4185
rect 1398 4111 1454 4120
rect 1398 3904 1454 3913
rect 1398 3839 1454 3848
rect 1412 3534 1440 3839
rect 1400 3528 1452 3534
rect 1400 3470 1452 3476
rect 1400 3392 1452 3398
rect 1400 3334 1452 3340
rect 1308 2440 1360 2446
rect 1308 2382 1360 2388
rect 848 2032 900 2038
rect 848 1974 900 1980
rect 1412 1057 1440 3334
rect 1504 2417 1532 5510
rect 1596 4026 1624 6054
rect 1688 4146 1716 8434
rect 1768 7812 1820 7818
rect 1768 7754 1820 7760
rect 1780 7177 1808 7754
rect 1766 7168 1822 7177
rect 1766 7103 1822 7112
rect 1768 6996 1820 7002
rect 1768 6938 1820 6944
rect 1780 4826 1808 6938
rect 1768 4820 1820 4826
rect 1768 4762 1820 4768
rect 1768 4684 1820 4690
rect 1768 4626 1820 4632
rect 1676 4140 1728 4146
rect 1676 4082 1728 4088
rect 1596 3998 1716 4026
rect 1688 2650 1716 3998
rect 1676 2644 1728 2650
rect 1676 2586 1728 2592
rect 1676 2440 1728 2446
rect 1490 2408 1546 2417
rect 1676 2382 1728 2388
rect 1490 2343 1546 2352
rect 1688 1698 1716 2382
rect 1780 2292 1808 4626
rect 1872 4214 1900 8774
rect 1950 8735 2006 8744
rect 2056 8294 2084 9030
rect 2134 8936 2190 8945
rect 2134 8871 2190 8880
rect 2228 8900 2280 8906
rect 2148 8634 2176 8871
rect 2228 8842 2280 8848
rect 2240 8673 2268 8842
rect 2226 8664 2282 8673
rect 2136 8628 2188 8634
rect 2226 8599 2228 8608
rect 2136 8570 2188 8576
rect 2280 8599 2282 8608
rect 2228 8570 2280 8576
rect 2240 8362 2268 8570
rect 2332 8514 2360 12396
rect 2516 11898 2544 12718
rect 2608 12209 2636 12838
rect 2594 12200 2650 12209
rect 2700 12170 2728 12922
rect 2962 12880 3018 12889
rect 2780 12844 2832 12850
rect 3068 12850 3096 14980
rect 3146 14920 3202 14929
rect 3146 14855 3202 14864
rect 3160 13530 3188 14855
rect 3252 14822 3280 15574
rect 3240 14816 3292 14822
rect 3240 14758 3292 14764
rect 3252 14074 3280 14758
rect 3240 14068 3292 14074
rect 3240 14010 3292 14016
rect 3240 13864 3292 13870
rect 3240 13806 3292 13812
rect 3148 13524 3200 13530
rect 3148 13466 3200 13472
rect 3148 13320 3200 13326
rect 3148 13262 3200 13268
rect 2962 12815 3018 12824
rect 3056 12844 3108 12850
rect 2780 12786 2832 12792
rect 2792 12753 2820 12786
rect 2976 12782 3004 12815
rect 3056 12786 3108 12792
rect 2964 12776 3016 12782
rect 2778 12744 2834 12753
rect 2964 12718 3016 12724
rect 2778 12679 2834 12688
rect 2870 12608 2926 12617
rect 2870 12543 2926 12552
rect 2594 12135 2650 12144
rect 2688 12164 2740 12170
rect 2688 12106 2740 12112
rect 2884 12084 2912 12543
rect 2884 12056 3004 12084
rect 2610 11996 2918 12005
rect 2610 11994 2616 11996
rect 2672 11994 2696 11996
rect 2752 11994 2776 11996
rect 2832 11994 2856 11996
rect 2912 11994 2918 11996
rect 2672 11942 2674 11994
rect 2854 11942 2856 11994
rect 2610 11940 2616 11942
rect 2672 11940 2696 11942
rect 2752 11940 2776 11942
rect 2832 11940 2856 11942
rect 2912 11940 2918 11942
rect 2610 11931 2918 11940
rect 2504 11892 2556 11898
rect 2504 11834 2556 11840
rect 2596 11620 2648 11626
rect 2596 11562 2648 11568
rect 2504 11552 2556 11558
rect 2504 11494 2556 11500
rect 2516 10826 2544 11494
rect 2608 11354 2636 11562
rect 2872 11552 2924 11558
rect 2872 11494 2924 11500
rect 2596 11348 2648 11354
rect 2596 11290 2648 11296
rect 2884 11132 2912 11494
rect 2976 11286 3004 12056
rect 3056 11756 3108 11762
rect 3056 11698 3108 11704
rect 2964 11280 3016 11286
rect 2964 11222 3016 11228
rect 2884 11104 3004 11132
rect 2610 10908 2918 10917
rect 2610 10906 2616 10908
rect 2672 10906 2696 10908
rect 2752 10906 2776 10908
rect 2832 10906 2856 10908
rect 2912 10906 2918 10908
rect 2672 10854 2674 10906
rect 2854 10854 2856 10906
rect 2610 10852 2616 10854
rect 2672 10852 2696 10854
rect 2752 10852 2776 10854
rect 2832 10852 2856 10854
rect 2912 10852 2918 10854
rect 2610 10843 2918 10852
rect 2424 10798 2544 10826
rect 2596 10804 2648 10810
rect 2424 9722 2452 10798
rect 2596 10746 2648 10752
rect 2502 10704 2558 10713
rect 2502 10639 2558 10648
rect 2412 9716 2464 9722
rect 2412 9658 2464 9664
rect 2410 9616 2466 9625
rect 2410 9551 2412 9560
rect 2464 9551 2466 9560
rect 2412 9522 2464 9528
rect 2424 9178 2452 9522
rect 2516 9178 2544 10639
rect 2608 10198 2636 10746
rect 2872 10736 2924 10742
rect 2872 10678 2924 10684
rect 2778 10432 2834 10441
rect 2778 10367 2834 10376
rect 2596 10192 2648 10198
rect 2596 10134 2648 10140
rect 2688 9988 2740 9994
rect 2792 9976 2820 10367
rect 2884 10130 2912 10678
rect 2872 10124 2924 10130
rect 2872 10066 2924 10072
rect 2740 9948 2820 9976
rect 2688 9930 2740 9936
rect 2610 9820 2918 9829
rect 2610 9818 2616 9820
rect 2672 9818 2696 9820
rect 2752 9818 2776 9820
rect 2832 9818 2856 9820
rect 2912 9818 2918 9820
rect 2672 9766 2674 9818
rect 2854 9766 2856 9818
rect 2610 9764 2616 9766
rect 2672 9764 2696 9766
rect 2752 9764 2776 9766
rect 2832 9764 2856 9766
rect 2912 9764 2918 9766
rect 2610 9755 2918 9764
rect 2596 9716 2648 9722
rect 2596 9658 2648 9664
rect 2608 9489 2636 9658
rect 2872 9648 2924 9654
rect 2870 9616 2872 9625
rect 2924 9616 2926 9625
rect 2780 9580 2832 9586
rect 2870 9551 2926 9560
rect 2976 9568 3004 11104
rect 3068 11082 3096 11698
rect 3056 11076 3108 11082
rect 3056 11018 3108 11024
rect 3054 10568 3110 10577
rect 3054 10503 3110 10512
rect 3068 10062 3096 10503
rect 3056 10056 3108 10062
rect 3056 9998 3108 10004
rect 3056 9580 3108 9586
rect 2976 9540 3056 9568
rect 2780 9522 2832 9528
rect 3056 9522 3108 9528
rect 2594 9480 2650 9489
rect 2594 9415 2650 9424
rect 2688 9376 2740 9382
rect 2688 9318 2740 9324
rect 2412 9172 2464 9178
rect 2412 9114 2464 9120
rect 2504 9172 2556 9178
rect 2504 9114 2556 9120
rect 2502 9072 2558 9081
rect 2502 9007 2558 9016
rect 2412 8900 2464 8906
rect 2412 8842 2464 8848
rect 2424 8634 2452 8842
rect 2412 8628 2464 8634
rect 2412 8570 2464 8576
rect 2332 8498 2452 8514
rect 2332 8492 2464 8498
rect 2332 8486 2412 8492
rect 2412 8434 2464 8440
rect 2320 8424 2372 8430
rect 2372 8372 2452 8378
rect 2320 8366 2452 8372
rect 2228 8356 2280 8362
rect 2332 8350 2452 8366
rect 2228 8298 2280 8304
rect 2044 8288 2096 8294
rect 2044 8230 2096 8236
rect 2320 8288 2372 8294
rect 2320 8230 2372 8236
rect 1950 8188 2258 8197
rect 1950 8186 1956 8188
rect 2012 8186 2036 8188
rect 2092 8186 2116 8188
rect 2172 8186 2196 8188
rect 2252 8186 2258 8188
rect 2012 8134 2014 8186
rect 2194 8134 2196 8186
rect 1950 8132 1956 8134
rect 2012 8132 2036 8134
rect 2092 8132 2116 8134
rect 2172 8132 2196 8134
rect 2252 8132 2258 8134
rect 1950 8123 2258 8132
rect 1950 7100 2258 7109
rect 1950 7098 1956 7100
rect 2012 7098 2036 7100
rect 2092 7098 2116 7100
rect 2172 7098 2196 7100
rect 2252 7098 2258 7100
rect 2012 7046 2014 7098
rect 2194 7046 2196 7098
rect 1950 7044 1956 7046
rect 2012 7044 2036 7046
rect 2092 7044 2116 7046
rect 2172 7044 2196 7046
rect 2252 7044 2258 7046
rect 1950 7035 2258 7044
rect 2332 6866 2360 8230
rect 2320 6860 2372 6866
rect 2320 6802 2372 6808
rect 2226 6760 2282 6769
rect 2226 6695 2282 6704
rect 2240 6225 2268 6695
rect 2226 6216 2282 6225
rect 2226 6151 2282 6160
rect 1950 6012 2258 6021
rect 1950 6010 1956 6012
rect 2012 6010 2036 6012
rect 2092 6010 2116 6012
rect 2172 6010 2196 6012
rect 2252 6010 2258 6012
rect 2012 5958 2014 6010
rect 2194 5958 2196 6010
rect 1950 5956 1956 5958
rect 2012 5956 2036 5958
rect 2092 5956 2116 5958
rect 2172 5956 2196 5958
rect 2252 5956 2258 5958
rect 1950 5947 2258 5956
rect 2332 5794 2360 6802
rect 2424 6769 2452 8350
rect 2516 7274 2544 9007
rect 2700 8838 2728 9318
rect 2792 8838 2820 9522
rect 2872 9512 2924 9518
rect 2872 9454 2924 9460
rect 2962 9480 3018 9489
rect 2688 8832 2740 8838
rect 2688 8774 2740 8780
rect 2780 8832 2832 8838
rect 2884 8820 2912 9454
rect 2962 9415 3018 9424
rect 2976 9160 3004 9415
rect 3068 9353 3096 9522
rect 3054 9344 3110 9353
rect 3054 9279 3110 9288
rect 2976 9132 3096 9160
rect 2962 9072 3018 9081
rect 2962 9007 3018 9016
rect 2976 8974 3004 9007
rect 2964 8968 3016 8974
rect 2964 8910 3016 8916
rect 2884 8792 3004 8820
rect 2780 8774 2832 8780
rect 2610 8732 2918 8741
rect 2610 8730 2616 8732
rect 2672 8730 2696 8732
rect 2752 8730 2776 8732
rect 2832 8730 2856 8732
rect 2912 8730 2918 8732
rect 2672 8678 2674 8730
rect 2854 8678 2856 8730
rect 2610 8676 2616 8678
rect 2672 8676 2696 8678
rect 2752 8676 2776 8678
rect 2832 8676 2856 8678
rect 2912 8676 2918 8678
rect 2610 8667 2918 8676
rect 2596 8628 2648 8634
rect 2648 8588 2820 8616
rect 2596 8570 2648 8576
rect 2594 8528 2650 8537
rect 2594 8463 2650 8472
rect 2608 8430 2636 8463
rect 2596 8424 2648 8430
rect 2596 8366 2648 8372
rect 2688 8288 2740 8294
rect 2688 8230 2740 8236
rect 2700 7834 2728 8230
rect 2792 8090 2820 8588
rect 2976 8514 3004 8792
rect 2884 8486 3004 8514
rect 2780 8084 2832 8090
rect 2780 8026 2832 8032
rect 2884 8022 2912 8486
rect 2964 8424 3016 8430
rect 3068 8412 3096 9132
rect 3016 8384 3096 8412
rect 2964 8366 3016 8372
rect 2872 8016 2924 8022
rect 2872 7958 2924 7964
rect 2700 7806 2820 7834
rect 2792 7750 2820 7806
rect 2780 7744 2832 7750
rect 2780 7686 2832 7692
rect 2610 7644 2918 7653
rect 2610 7642 2616 7644
rect 2672 7642 2696 7644
rect 2752 7642 2776 7644
rect 2832 7642 2856 7644
rect 2912 7642 2918 7644
rect 2672 7590 2674 7642
rect 2854 7590 2856 7642
rect 2610 7588 2616 7590
rect 2672 7588 2696 7590
rect 2752 7588 2776 7590
rect 2832 7588 2856 7590
rect 2912 7588 2918 7590
rect 2610 7579 2918 7588
rect 2504 7268 2556 7274
rect 2504 7210 2556 7216
rect 2504 6996 2556 7002
rect 2504 6938 2556 6944
rect 2410 6760 2466 6769
rect 2410 6695 2466 6704
rect 2516 5914 2544 6938
rect 2610 6556 2918 6565
rect 2610 6554 2616 6556
rect 2672 6554 2696 6556
rect 2752 6554 2776 6556
rect 2832 6554 2856 6556
rect 2912 6554 2918 6556
rect 2672 6502 2674 6554
rect 2854 6502 2856 6554
rect 2610 6500 2616 6502
rect 2672 6500 2696 6502
rect 2752 6500 2776 6502
rect 2832 6500 2856 6502
rect 2912 6500 2918 6502
rect 2610 6491 2918 6500
rect 2872 6384 2924 6390
rect 2872 6326 2924 6332
rect 2596 6180 2648 6186
rect 2596 6122 2648 6128
rect 2504 5908 2556 5914
rect 2504 5850 2556 5856
rect 2608 5896 2636 6122
rect 2688 5908 2740 5914
rect 2608 5868 2688 5896
rect 2332 5766 2544 5794
rect 2412 5704 2464 5710
rect 2412 5646 2464 5652
rect 2320 5636 2372 5642
rect 2320 5578 2372 5584
rect 1950 4924 2258 4933
rect 1950 4922 1956 4924
rect 2012 4922 2036 4924
rect 2092 4922 2116 4924
rect 2172 4922 2196 4924
rect 2252 4922 2258 4924
rect 2012 4870 2014 4922
rect 2194 4870 2196 4922
rect 1950 4868 1956 4870
rect 2012 4868 2036 4870
rect 2092 4868 2116 4870
rect 2172 4868 2196 4870
rect 2252 4868 2258 4870
rect 1950 4859 2258 4868
rect 1952 4820 2004 4826
rect 1952 4762 2004 4768
rect 1860 4208 1912 4214
rect 1860 4150 1912 4156
rect 1964 4026 1992 4762
rect 2228 4140 2280 4146
rect 2332 4128 2360 5578
rect 2424 5302 2452 5646
rect 2412 5296 2464 5302
rect 2412 5238 2464 5244
rect 2516 4826 2544 5766
rect 2608 5710 2636 5868
rect 2688 5850 2740 5856
rect 2884 5778 2912 6326
rect 2872 5772 2924 5778
rect 2872 5714 2924 5720
rect 2596 5704 2648 5710
rect 2596 5646 2648 5652
rect 2610 5468 2918 5477
rect 2610 5466 2616 5468
rect 2672 5466 2696 5468
rect 2752 5466 2776 5468
rect 2832 5466 2856 5468
rect 2912 5466 2918 5468
rect 2672 5414 2674 5466
rect 2854 5414 2856 5466
rect 2610 5412 2616 5414
rect 2672 5412 2696 5414
rect 2752 5412 2776 5414
rect 2832 5412 2856 5414
rect 2912 5412 2918 5414
rect 2610 5403 2918 5412
rect 2778 4856 2834 4865
rect 2504 4820 2556 4826
rect 2778 4791 2834 4800
rect 2504 4762 2556 4768
rect 2792 4758 2820 4791
rect 2780 4752 2832 4758
rect 2780 4694 2832 4700
rect 2412 4616 2464 4622
rect 2412 4558 2464 4564
rect 2280 4100 2360 4128
rect 2228 4082 2280 4088
rect 1872 3998 1992 4026
rect 2320 4004 2372 4010
rect 1872 3720 1900 3998
rect 2320 3946 2372 3952
rect 1950 3836 2258 3845
rect 1950 3834 1956 3836
rect 2012 3834 2036 3836
rect 2092 3834 2116 3836
rect 2172 3834 2196 3836
rect 2252 3834 2258 3836
rect 2012 3782 2014 3834
rect 2194 3782 2196 3834
rect 1950 3780 1956 3782
rect 2012 3780 2036 3782
rect 2092 3780 2116 3782
rect 2172 3780 2196 3782
rect 2252 3780 2258 3782
rect 1950 3771 2258 3780
rect 1872 3692 1992 3720
rect 1860 3528 1912 3534
rect 1860 3470 1912 3476
rect 1872 2446 1900 3470
rect 1964 3398 1992 3692
rect 2332 3670 2360 3946
rect 2424 3913 2452 4558
rect 2610 4380 2918 4389
rect 2610 4378 2616 4380
rect 2672 4378 2696 4380
rect 2752 4378 2776 4380
rect 2832 4378 2856 4380
rect 2912 4378 2918 4380
rect 2672 4326 2674 4378
rect 2854 4326 2856 4378
rect 2610 4324 2616 4326
rect 2672 4324 2696 4326
rect 2752 4324 2776 4326
rect 2832 4324 2856 4326
rect 2912 4324 2918 4326
rect 2610 4315 2918 4324
rect 2596 4276 2648 4282
rect 2516 4236 2596 4264
rect 2410 3904 2466 3913
rect 2410 3839 2466 3848
rect 2320 3664 2372 3670
rect 2320 3606 2372 3612
rect 1952 3392 2004 3398
rect 1952 3334 2004 3340
rect 2412 3052 2464 3058
rect 2412 2994 2464 3000
rect 1950 2748 2258 2757
rect 1950 2746 1956 2748
rect 2012 2746 2036 2748
rect 2092 2746 2116 2748
rect 2172 2746 2196 2748
rect 2252 2746 2258 2748
rect 2012 2694 2014 2746
rect 2194 2694 2196 2746
rect 1950 2692 1956 2694
rect 2012 2692 2036 2694
rect 2092 2692 2116 2694
rect 2172 2692 2196 2694
rect 2252 2692 2258 2694
rect 1950 2683 2258 2692
rect 2424 2530 2452 2994
rect 2516 2990 2544 4236
rect 2596 4218 2648 4224
rect 2976 3942 3004 8366
rect 3056 8288 3108 8294
rect 3056 8230 3108 8236
rect 3068 8129 3096 8230
rect 3054 8120 3110 8129
rect 3054 8055 3110 8064
rect 3056 7744 3108 7750
rect 3056 7686 3108 7692
rect 3068 5370 3096 7686
rect 3160 7002 3188 13262
rect 3252 13025 3280 13806
rect 3238 13016 3294 13025
rect 3238 12951 3294 12960
rect 3252 12850 3280 12951
rect 3344 12889 3372 18430
rect 3608 18012 3660 18018
rect 3608 17954 3660 17960
rect 3516 17536 3568 17542
rect 3516 17478 3568 17484
rect 3424 14000 3476 14006
rect 3424 13942 3476 13948
rect 3330 12880 3386 12889
rect 3240 12844 3292 12850
rect 3330 12815 3386 12824
rect 3240 12786 3292 12792
rect 3240 12640 3292 12646
rect 3240 12582 3292 12588
rect 3148 6996 3200 7002
rect 3148 6938 3200 6944
rect 3148 6724 3200 6730
rect 3148 6666 3200 6672
rect 3160 6390 3188 6666
rect 3148 6384 3200 6390
rect 3148 6326 3200 6332
rect 3148 6248 3200 6254
rect 3148 6190 3200 6196
rect 3056 5364 3108 5370
rect 3056 5306 3108 5312
rect 3054 5264 3110 5273
rect 3054 5199 3056 5208
rect 3108 5199 3110 5208
rect 3056 5170 3108 5176
rect 2964 3936 3016 3942
rect 2964 3878 3016 3884
rect 3068 3754 3096 5170
rect 2884 3726 3096 3754
rect 2884 3602 2912 3726
rect 3056 3664 3108 3670
rect 2976 3612 3056 3618
rect 2976 3606 3108 3612
rect 2872 3596 2924 3602
rect 2872 3538 2924 3544
rect 2976 3590 3096 3606
rect 2688 3528 2740 3534
rect 2976 3482 3004 3590
rect 3056 3528 3108 3534
rect 2740 3476 3004 3482
rect 2688 3470 3004 3476
rect 2700 3454 3004 3470
rect 3054 3496 3056 3505
rect 3108 3496 3110 3505
rect 3054 3431 3110 3440
rect 2964 3392 3016 3398
rect 2964 3334 3016 3340
rect 2610 3292 2918 3301
rect 2610 3290 2616 3292
rect 2672 3290 2696 3292
rect 2752 3290 2776 3292
rect 2832 3290 2856 3292
rect 2912 3290 2918 3292
rect 2672 3238 2674 3290
rect 2854 3238 2856 3290
rect 2610 3236 2616 3238
rect 2672 3236 2696 3238
rect 2752 3236 2776 3238
rect 2832 3236 2856 3238
rect 2912 3236 2918 3238
rect 2610 3227 2918 3236
rect 2778 3088 2834 3097
rect 2976 3058 3004 3334
rect 3160 3062 3188 6190
rect 3252 4690 3280 12582
rect 3436 12481 3464 13942
rect 3528 12918 3556 17478
rect 3620 15434 3648 17954
rect 3712 17270 3740 19200
rect 5816 18828 5868 18834
rect 5816 18770 5868 18776
rect 5632 18556 5684 18562
rect 5632 18498 5684 18504
rect 5264 18352 5316 18358
rect 5264 18294 5316 18300
rect 4250 17912 4306 17921
rect 4250 17847 4306 17856
rect 3976 17672 4028 17678
rect 3976 17614 4028 17620
rect 3882 17368 3938 17377
rect 3882 17303 3938 17312
rect 3700 17264 3752 17270
rect 3700 17206 3752 17212
rect 3698 16280 3754 16289
rect 3698 16215 3754 16224
rect 3608 15428 3660 15434
rect 3608 15370 3660 15376
rect 3608 14340 3660 14346
rect 3608 14282 3660 14288
rect 3620 13734 3648 14282
rect 3608 13728 3660 13734
rect 3608 13670 3660 13676
rect 3516 12912 3568 12918
rect 3516 12854 3568 12860
rect 3422 12472 3478 12481
rect 3422 12407 3478 12416
rect 3528 12186 3556 12854
rect 3608 12640 3660 12646
rect 3608 12582 3660 12588
rect 3332 12164 3384 12170
rect 3332 12106 3384 12112
rect 3436 12158 3556 12186
rect 3344 9761 3372 12106
rect 3436 11830 3464 12158
rect 3516 12096 3568 12102
rect 3516 12038 3568 12044
rect 3424 11824 3476 11830
rect 3424 11766 3476 11772
rect 3436 11014 3464 11766
rect 3528 11694 3556 12038
rect 3620 11937 3648 12582
rect 3712 12306 3740 16215
rect 3896 15570 3924 17303
rect 3884 15564 3936 15570
rect 3884 15506 3936 15512
rect 3884 14952 3936 14958
rect 3884 14894 3936 14900
rect 3896 13938 3924 14894
rect 3988 14890 4016 17614
rect 4160 15972 4212 15978
rect 4160 15914 4212 15920
rect 4066 15600 4122 15609
rect 4066 15535 4068 15544
rect 4120 15535 4122 15544
rect 4068 15506 4120 15512
rect 4172 15502 4200 15914
rect 4160 15496 4212 15502
rect 4066 15464 4122 15473
rect 4160 15438 4212 15444
rect 4066 15399 4122 15408
rect 3976 14884 4028 14890
rect 3976 14826 4028 14832
rect 3884 13932 3936 13938
rect 3884 13874 3936 13880
rect 3792 13252 3844 13258
rect 3792 13194 3844 13200
rect 3804 12442 3832 13194
rect 3896 12646 3924 13874
rect 3976 13728 4028 13734
rect 3976 13670 4028 13676
rect 3884 12640 3936 12646
rect 3884 12582 3936 12588
rect 3882 12472 3938 12481
rect 3792 12436 3844 12442
rect 3882 12407 3938 12416
rect 3792 12378 3844 12384
rect 3700 12300 3752 12306
rect 3700 12242 3752 12248
rect 3700 12164 3752 12170
rect 3700 12106 3752 12112
rect 3606 11928 3662 11937
rect 3606 11863 3662 11872
rect 3608 11756 3660 11762
rect 3608 11698 3660 11704
rect 3516 11688 3568 11694
rect 3516 11630 3568 11636
rect 3424 11008 3476 11014
rect 3424 10950 3476 10956
rect 3514 10976 3570 10985
rect 3514 10911 3570 10920
rect 3424 10804 3476 10810
rect 3424 10746 3476 10752
rect 3330 9752 3386 9761
rect 3330 9687 3386 9696
rect 3332 9512 3384 9518
rect 3332 9454 3384 9460
rect 3344 9353 3372 9454
rect 3330 9344 3386 9353
rect 3330 9279 3386 9288
rect 3436 9178 3464 10746
rect 3528 10470 3556 10911
rect 3620 10810 3648 11698
rect 3712 11354 3740 12106
rect 3790 12064 3846 12073
rect 3790 11999 3846 12008
rect 3700 11348 3752 11354
rect 3700 11290 3752 11296
rect 3608 10804 3660 10810
rect 3608 10746 3660 10752
rect 3608 10668 3660 10674
rect 3608 10610 3660 10616
rect 3516 10464 3568 10470
rect 3516 10406 3568 10412
rect 3528 10169 3556 10406
rect 3514 10160 3570 10169
rect 3514 10095 3570 10104
rect 3620 10062 3648 10610
rect 3700 10464 3752 10470
rect 3700 10406 3752 10412
rect 3608 10056 3660 10062
rect 3606 10024 3608 10033
rect 3660 10024 3662 10033
rect 3606 9959 3662 9968
rect 3516 9920 3568 9926
rect 3514 9888 3516 9897
rect 3568 9888 3570 9897
rect 3514 9823 3570 9832
rect 3516 9512 3568 9518
rect 3516 9454 3568 9460
rect 3606 9480 3662 9489
rect 3424 9172 3476 9178
rect 3344 9132 3424 9160
rect 3344 6730 3372 9132
rect 3424 9114 3476 9120
rect 3422 8800 3478 8809
rect 3422 8735 3478 8744
rect 3436 8566 3464 8735
rect 3528 8650 3556 9454
rect 3606 9415 3662 9424
rect 3620 9382 3648 9415
rect 3608 9376 3660 9382
rect 3608 9318 3660 9324
rect 3608 8900 3660 8906
rect 3608 8842 3660 8848
rect 3620 8809 3648 8842
rect 3606 8800 3662 8809
rect 3606 8735 3662 8744
rect 3528 8622 3648 8650
rect 3424 8560 3476 8566
rect 3424 8502 3476 8508
rect 3514 8528 3570 8537
rect 3514 8463 3516 8472
rect 3568 8463 3570 8472
rect 3516 8434 3568 8440
rect 3514 8392 3570 8401
rect 3514 8327 3570 8336
rect 3424 6996 3476 7002
rect 3424 6938 3476 6944
rect 3332 6724 3384 6730
rect 3332 6666 3384 6672
rect 3330 6488 3386 6497
rect 3330 6423 3386 6432
rect 3344 6390 3372 6423
rect 3332 6384 3384 6390
rect 3332 6326 3384 6332
rect 3332 5908 3384 5914
rect 3332 5850 3384 5856
rect 3240 4684 3292 4690
rect 3240 4626 3292 4632
rect 3344 4570 3372 5850
rect 3436 5778 3464 6938
rect 3528 6390 3556 8327
rect 3620 8129 3648 8622
rect 3606 8120 3662 8129
rect 3606 8055 3662 8064
rect 3608 7948 3660 7954
rect 3608 7890 3660 7896
rect 3620 6866 3648 7890
rect 3608 6860 3660 6866
rect 3608 6802 3660 6808
rect 3712 6712 3740 10406
rect 3804 9654 3832 11999
rect 3896 11830 3924 12407
rect 3884 11824 3936 11830
rect 3884 11766 3936 11772
rect 3884 11144 3936 11150
rect 3884 11086 3936 11092
rect 3896 10198 3924 11086
rect 3988 10674 4016 13670
rect 4080 13569 4108 15399
rect 4066 13560 4122 13569
rect 4066 13495 4122 13504
rect 4068 13320 4120 13326
rect 4068 13262 4120 13268
rect 4080 11898 4108 13262
rect 4264 13258 4292 17847
rect 4436 17808 4488 17814
rect 4436 17750 4488 17756
rect 4344 15496 4396 15502
rect 4344 15438 4396 15444
rect 4252 13252 4304 13258
rect 4252 13194 4304 13200
rect 4250 13152 4306 13161
rect 4250 13087 4306 13096
rect 4264 12458 4292 13087
rect 4356 12617 4384 15438
rect 4448 14657 4476 17750
rect 4804 17740 4856 17746
rect 4804 17682 4856 17688
rect 4620 16244 4672 16250
rect 4620 16186 4672 16192
rect 4632 15026 4660 16186
rect 4710 16144 4766 16153
rect 4710 16079 4766 16088
rect 4724 15570 4752 16079
rect 4712 15564 4764 15570
rect 4712 15506 4764 15512
rect 4528 15020 4580 15026
rect 4528 14962 4580 14968
rect 4620 15020 4672 15026
rect 4620 14962 4672 14968
rect 4434 14648 4490 14657
rect 4434 14583 4490 14592
rect 4434 14512 4490 14521
rect 4434 14447 4490 14456
rect 4342 12608 4398 12617
rect 4342 12543 4398 12552
rect 4160 12436 4212 12442
rect 4264 12430 4384 12458
rect 4160 12378 4212 12384
rect 4068 11892 4120 11898
rect 4068 11834 4120 11840
rect 4066 11792 4122 11801
rect 4172 11762 4200 12378
rect 4252 12232 4304 12238
rect 4252 12174 4304 12180
rect 4264 11801 4292 12174
rect 4250 11792 4306 11801
rect 4066 11727 4122 11736
rect 4160 11756 4212 11762
rect 4080 11286 4108 11727
rect 4250 11727 4306 11736
rect 4160 11698 4212 11704
rect 4252 11688 4304 11694
rect 4252 11630 4304 11636
rect 4160 11348 4212 11354
rect 4160 11290 4212 11296
rect 4068 11280 4120 11286
rect 4068 11222 4120 11228
rect 3976 10668 4028 10674
rect 3976 10610 4028 10616
rect 3976 10532 4028 10538
rect 4028 10492 4108 10520
rect 3976 10474 4028 10480
rect 3974 10432 4030 10441
rect 3974 10367 4030 10376
rect 3988 10266 4016 10367
rect 3976 10260 4028 10266
rect 3976 10202 4028 10208
rect 3884 10192 3936 10198
rect 3884 10134 3936 10140
rect 3974 10160 4030 10169
rect 3792 9648 3844 9654
rect 3792 9590 3844 9596
rect 3896 9586 3924 10134
rect 3974 10095 4030 10104
rect 3884 9580 3936 9586
rect 3884 9522 3936 9528
rect 3882 9344 3938 9353
rect 3882 9279 3938 9288
rect 3792 9172 3844 9178
rect 3792 9114 3844 9120
rect 3804 7857 3832 9114
rect 3896 9110 3924 9279
rect 3884 9104 3936 9110
rect 3884 9046 3936 9052
rect 3884 8900 3936 8906
rect 3884 8842 3936 8848
rect 3896 8634 3924 8842
rect 3884 8628 3936 8634
rect 3884 8570 3936 8576
rect 3882 8528 3938 8537
rect 3882 8463 3938 8472
rect 3896 8430 3924 8463
rect 3884 8424 3936 8430
rect 3884 8366 3936 8372
rect 3988 8276 4016 10095
rect 4080 9353 4108 10492
rect 4066 9344 4122 9353
rect 4066 9279 4122 9288
rect 4172 9178 4200 11290
rect 4264 10690 4292 11630
rect 4356 10810 4384 12430
rect 4448 12238 4476 14447
rect 4540 14385 4568 14962
rect 4712 14408 4764 14414
rect 4526 14376 4582 14385
rect 4712 14350 4764 14356
rect 4526 14311 4582 14320
rect 4620 14068 4672 14074
rect 4620 14010 4672 14016
rect 4528 13320 4580 13326
rect 4528 13262 4580 13268
rect 4436 12232 4488 12238
rect 4436 12174 4488 12180
rect 4436 11756 4488 11762
rect 4436 11698 4488 11704
rect 4448 11393 4476 11698
rect 4434 11384 4490 11393
rect 4434 11319 4490 11328
rect 4436 11280 4488 11286
rect 4436 11222 4488 11228
rect 4448 10996 4476 11222
rect 4540 11064 4568 13262
rect 4632 12850 4660 14010
rect 4724 13841 4752 14350
rect 4816 14090 4844 17682
rect 4896 16992 4948 16998
rect 4896 16934 4948 16940
rect 4908 15502 4936 16934
rect 4988 16720 5040 16726
rect 4988 16662 5040 16668
rect 4896 15496 4948 15502
rect 4896 15438 4948 15444
rect 4894 15192 4950 15201
rect 4894 15127 4950 15136
rect 4908 14278 4936 15127
rect 5000 14414 5028 16662
rect 5172 16244 5224 16250
rect 5172 16186 5224 16192
rect 5184 15502 5212 16186
rect 5172 15496 5224 15502
rect 5092 15456 5172 15484
rect 4988 14408 5040 14414
rect 4988 14350 5040 14356
rect 4896 14272 4948 14278
rect 4894 14240 4896 14249
rect 4948 14240 4950 14249
rect 4894 14175 4950 14184
rect 4816 14062 4936 14090
rect 4804 13932 4856 13938
rect 4804 13874 4856 13880
rect 4710 13832 4766 13841
rect 4710 13767 4766 13776
rect 4712 13524 4764 13530
rect 4712 13466 4764 13472
rect 4724 12918 4752 13466
rect 4712 12912 4764 12918
rect 4712 12854 4764 12860
rect 4620 12844 4672 12850
rect 4620 12786 4672 12792
rect 4620 12708 4672 12714
rect 4620 12650 4672 12656
rect 4632 12481 4660 12650
rect 4618 12472 4674 12481
rect 4618 12407 4674 12416
rect 4618 12336 4674 12345
rect 4618 12271 4674 12280
rect 4632 11354 4660 12271
rect 4724 11558 4752 12854
rect 4816 11801 4844 13874
rect 4802 11792 4858 11801
rect 4802 11727 4858 11736
rect 4712 11552 4764 11558
rect 4712 11494 4764 11500
rect 4710 11384 4766 11393
rect 4620 11348 4672 11354
rect 4710 11319 4766 11328
rect 4620 11290 4672 11296
rect 4618 11248 4674 11257
rect 4618 11183 4620 11192
rect 4672 11183 4674 11192
rect 4620 11154 4672 11160
rect 4540 11036 4660 11064
rect 4448 10968 4568 10996
rect 4344 10804 4396 10810
rect 4344 10746 4396 10752
rect 4540 10724 4568 10968
rect 4448 10696 4568 10724
rect 4264 10674 4384 10690
rect 4264 10668 4396 10674
rect 4264 10662 4344 10668
rect 4344 10610 4396 10616
rect 4252 10600 4304 10606
rect 4252 10542 4304 10548
rect 4264 10062 4292 10542
rect 4344 10260 4396 10266
rect 4344 10202 4396 10208
rect 4252 10056 4304 10062
rect 4356 10033 4384 10202
rect 4252 9998 4304 10004
rect 4342 10024 4398 10033
rect 4264 9722 4292 9998
rect 4342 9959 4398 9968
rect 4342 9752 4398 9761
rect 4252 9716 4304 9722
rect 4342 9687 4398 9696
rect 4252 9658 4304 9664
rect 4252 9512 4304 9518
rect 4252 9454 4304 9460
rect 4160 9172 4212 9178
rect 4160 9114 4212 9120
rect 4264 8974 4292 9454
rect 4068 8968 4120 8974
rect 4160 8968 4212 8974
rect 4068 8910 4120 8916
rect 4158 8936 4160 8945
rect 4252 8968 4304 8974
rect 4212 8936 4214 8945
rect 3896 8248 4016 8276
rect 3896 7954 3924 8248
rect 3974 8120 4030 8129
rect 3974 8055 4030 8064
rect 3884 7948 3936 7954
rect 3884 7890 3936 7896
rect 3790 7848 3846 7857
rect 3790 7783 3846 7792
rect 3884 7812 3936 7818
rect 3804 6798 3832 7783
rect 3884 7754 3936 7760
rect 3896 7041 3924 7754
rect 3988 7449 4016 8055
rect 3974 7440 4030 7449
rect 3974 7375 4030 7384
rect 3976 7200 4028 7206
rect 3976 7142 4028 7148
rect 3882 7032 3938 7041
rect 3882 6967 3938 6976
rect 3884 6928 3936 6934
rect 3884 6870 3936 6876
rect 3792 6792 3844 6798
rect 3792 6734 3844 6740
rect 3620 6684 3740 6712
rect 3620 6440 3648 6684
rect 3792 6656 3844 6662
rect 3792 6598 3844 6604
rect 3620 6412 3740 6440
rect 3516 6384 3568 6390
rect 3516 6326 3568 6332
rect 3608 6316 3660 6322
rect 3608 6258 3660 6264
rect 3514 6216 3570 6225
rect 3514 6151 3570 6160
rect 3528 6118 3556 6151
rect 3516 6112 3568 6118
rect 3516 6054 3568 6060
rect 3620 5914 3648 6258
rect 3608 5908 3660 5914
rect 3608 5850 3660 5856
rect 3424 5772 3476 5778
rect 3424 5714 3476 5720
rect 3608 5568 3660 5574
rect 3514 5536 3570 5545
rect 3608 5510 3660 5516
rect 3514 5471 3570 5480
rect 3424 5296 3476 5302
rect 3424 5238 3476 5244
rect 3252 4542 3372 4570
rect 3252 3466 3280 4542
rect 3330 4312 3386 4321
rect 3330 4247 3386 4256
rect 3240 3460 3292 3466
rect 3240 3402 3292 3408
rect 2778 3023 2780 3032
rect 2832 3023 2834 3032
rect 2964 3052 3016 3058
rect 2780 2994 2832 3000
rect 2964 2994 3016 3000
rect 3068 3034 3188 3062
rect 3344 3058 3372 4247
rect 3436 3369 3464 5238
rect 3422 3360 3478 3369
rect 3422 3295 3478 3304
rect 3332 3052 3384 3058
rect 2504 2984 2556 2990
rect 2504 2926 2556 2932
rect 2964 2848 3016 2854
rect 2964 2790 3016 2796
rect 2332 2502 2452 2530
rect 1860 2440 1912 2446
rect 1860 2382 1912 2388
rect 2044 2440 2096 2446
rect 2044 2382 2096 2388
rect 2056 2292 2084 2382
rect 1780 2264 2084 2292
rect 1676 1692 1728 1698
rect 1676 1634 1728 1640
rect 2332 1358 2360 2502
rect 2412 2440 2464 2446
rect 2412 2382 2464 2388
rect 2424 1465 2452 2382
rect 2504 2304 2556 2310
rect 2504 2246 2556 2252
rect 2410 1456 2466 1465
rect 2516 1442 2544 2246
rect 2610 2204 2918 2213
rect 2610 2202 2616 2204
rect 2672 2202 2696 2204
rect 2752 2202 2776 2204
rect 2832 2202 2856 2204
rect 2912 2202 2918 2204
rect 2672 2150 2674 2202
rect 2854 2150 2856 2202
rect 2610 2148 2616 2150
rect 2672 2148 2696 2150
rect 2752 2148 2776 2150
rect 2832 2148 2856 2150
rect 2912 2148 2918 2150
rect 2610 2139 2918 2148
rect 2594 1456 2650 1465
rect 2516 1414 2594 1442
rect 2410 1391 2466 1400
rect 2594 1391 2650 1400
rect 2320 1352 2372 1358
rect 2320 1294 2372 1300
rect 2976 1086 3004 2790
rect 3068 1834 3096 3034
rect 3332 2994 3384 3000
rect 3148 2984 3200 2990
rect 3148 2926 3200 2932
rect 3240 2984 3292 2990
rect 3240 2926 3292 2932
rect 3056 1828 3108 1834
rect 3056 1770 3108 1776
rect 2964 1080 3016 1086
rect 1398 1048 1454 1057
rect 2964 1022 3016 1028
rect 1398 983 1454 992
rect 3160 950 3188 2926
rect 3252 2145 3280 2926
rect 3436 2650 3464 3295
rect 3528 3058 3556 5471
rect 3620 5302 3648 5510
rect 3608 5296 3660 5302
rect 3608 5238 3660 5244
rect 3712 3194 3740 6412
rect 3700 3188 3752 3194
rect 3700 3130 3752 3136
rect 3516 3052 3568 3058
rect 3516 2994 3568 3000
rect 3804 2650 3832 6598
rect 3896 6066 3924 6870
rect 3988 6322 4016 7142
rect 4080 7002 4108 8910
rect 4252 8910 4304 8916
rect 4158 8871 4214 8880
rect 4160 8832 4212 8838
rect 4160 8774 4212 8780
rect 4252 8832 4304 8838
rect 4252 8774 4304 8780
rect 4068 6996 4120 7002
rect 4068 6938 4120 6944
rect 4066 6896 4122 6905
rect 4066 6831 4122 6840
rect 4080 6798 4108 6831
rect 4068 6792 4120 6798
rect 4068 6734 4120 6740
rect 4172 6440 4200 8774
rect 4264 8634 4292 8774
rect 4252 8628 4304 8634
rect 4252 8570 4304 8576
rect 4252 8492 4304 8498
rect 4356 8480 4384 9687
rect 4304 8452 4384 8480
rect 4252 8434 4304 8440
rect 4264 7290 4292 8434
rect 4344 8356 4396 8362
rect 4344 8298 4396 8304
rect 4356 7818 4384 8298
rect 4344 7812 4396 7818
rect 4344 7754 4396 7760
rect 4356 7410 4384 7754
rect 4344 7404 4396 7410
rect 4344 7346 4396 7352
rect 4264 7262 4384 7290
rect 4356 7002 4384 7262
rect 4344 6996 4396 7002
rect 4344 6938 4396 6944
rect 4344 6860 4396 6866
rect 4344 6802 4396 6808
rect 4252 6452 4304 6458
rect 4172 6412 4252 6440
rect 4252 6394 4304 6400
rect 4158 6352 4214 6361
rect 3976 6316 4028 6322
rect 4028 6276 4108 6304
rect 4158 6287 4214 6296
rect 3976 6258 4028 6264
rect 3974 6216 4030 6225
rect 3974 6151 3976 6160
rect 4028 6151 4030 6160
rect 3976 6122 4028 6128
rect 3896 6038 4016 6066
rect 3882 5808 3938 5817
rect 3882 5743 3938 5752
rect 3896 4282 3924 5743
rect 3988 5409 4016 6038
rect 4080 5953 4108 6276
rect 4066 5944 4122 5953
rect 4066 5879 4122 5888
rect 4068 5772 4120 5778
rect 4172 5760 4200 6287
rect 4120 5732 4200 5760
rect 4068 5714 4120 5720
rect 4160 5568 4212 5574
rect 4160 5510 4212 5516
rect 3974 5400 4030 5409
rect 3974 5335 4030 5344
rect 3988 5234 4016 5335
rect 4172 5234 4200 5510
rect 4356 5234 4384 6802
rect 4448 6798 4476 10696
rect 4632 10554 4660 11036
rect 4724 10742 4752 11319
rect 4908 11200 4936 14062
rect 4988 13796 5040 13802
rect 4988 13738 5040 13744
rect 5000 13530 5028 13738
rect 4988 13524 5040 13530
rect 4988 13466 5040 13472
rect 4986 13424 5042 13433
rect 4986 13359 5042 13368
rect 5000 12918 5028 13359
rect 4988 12912 5040 12918
rect 4988 12854 5040 12860
rect 4988 12232 5040 12238
rect 4988 12174 5040 12180
rect 4816 11172 4936 11200
rect 4816 11082 4844 11172
rect 4804 11076 4856 11082
rect 4804 11018 4856 11024
rect 5000 10810 5028 12174
rect 5092 11393 5120 15456
rect 5172 15438 5224 15444
rect 5276 15094 5304 18294
rect 5354 17232 5410 17241
rect 5354 17167 5410 17176
rect 5448 17196 5500 17202
rect 5368 17134 5396 17167
rect 5448 17138 5500 17144
rect 5356 17128 5408 17134
rect 5356 17070 5408 17076
rect 5460 16833 5488 17138
rect 5446 16824 5502 16833
rect 5446 16759 5502 16768
rect 5448 16652 5500 16658
rect 5448 16594 5500 16600
rect 5460 15706 5488 16594
rect 5356 15700 5408 15706
rect 5356 15642 5408 15648
rect 5448 15700 5500 15706
rect 5448 15642 5500 15648
rect 5368 15484 5396 15642
rect 5368 15456 5580 15484
rect 5552 15366 5580 15456
rect 5448 15360 5500 15366
rect 5448 15302 5500 15308
rect 5540 15360 5592 15366
rect 5540 15302 5592 15308
rect 5264 15088 5316 15094
rect 5460 15065 5488 15302
rect 5264 15030 5316 15036
rect 5446 15056 5502 15065
rect 5644 15008 5672 18498
rect 5828 18057 5856 18770
rect 6092 18760 6144 18766
rect 6092 18702 6144 18708
rect 5814 18048 5870 18057
rect 5814 17983 5870 17992
rect 5724 15700 5776 15706
rect 5724 15642 5776 15648
rect 5446 14991 5502 15000
rect 5552 14980 5672 15008
rect 5172 14408 5224 14414
rect 5172 14350 5224 14356
rect 5264 14408 5316 14414
rect 5264 14350 5316 14356
rect 5184 13870 5212 14350
rect 5172 13864 5224 13870
rect 5172 13806 5224 13812
rect 5172 13728 5224 13734
rect 5172 13670 5224 13676
rect 5184 13394 5212 13670
rect 5172 13388 5224 13394
rect 5172 13330 5224 13336
rect 5276 12434 5304 14350
rect 5354 14104 5410 14113
rect 5354 14039 5410 14048
rect 5368 14006 5396 14039
rect 5356 14000 5408 14006
rect 5356 13942 5408 13948
rect 5446 13968 5502 13977
rect 5446 13903 5502 13912
rect 5356 13864 5408 13870
rect 5356 13806 5408 13812
rect 5368 13530 5396 13806
rect 5460 13530 5488 13903
rect 5552 13870 5580 14980
rect 5632 14884 5684 14890
rect 5632 14826 5684 14832
rect 5540 13864 5592 13870
rect 5540 13806 5592 13812
rect 5538 13560 5594 13569
rect 5356 13524 5408 13530
rect 5356 13466 5408 13472
rect 5448 13524 5500 13530
rect 5538 13495 5594 13504
rect 5448 13466 5500 13472
rect 5552 13410 5580 13495
rect 5460 13394 5580 13410
rect 5448 13388 5580 13394
rect 5500 13382 5580 13388
rect 5448 13330 5500 13336
rect 5356 13252 5408 13258
rect 5356 13194 5408 13200
rect 5368 12850 5396 13194
rect 5644 13025 5672 14826
rect 5736 13938 5764 15642
rect 6000 14476 6052 14482
rect 6000 14418 6052 14424
rect 5908 14272 5960 14278
rect 5908 14214 5960 14220
rect 5920 13938 5948 14214
rect 5724 13932 5776 13938
rect 5724 13874 5776 13880
rect 5908 13932 5960 13938
rect 5908 13874 5960 13880
rect 5816 13864 5868 13870
rect 5816 13806 5868 13812
rect 5906 13832 5962 13841
rect 5724 13728 5776 13734
rect 5724 13670 5776 13676
rect 5630 13016 5686 13025
rect 5630 12951 5686 12960
rect 5356 12844 5408 12850
rect 5356 12786 5408 12792
rect 5448 12844 5500 12850
rect 5448 12786 5500 12792
rect 5632 12844 5684 12850
rect 5632 12786 5684 12792
rect 5276 12406 5396 12434
rect 5264 11892 5316 11898
rect 5264 11834 5316 11840
rect 5172 11756 5224 11762
rect 5172 11698 5224 11704
rect 5078 11384 5134 11393
rect 5078 11319 5134 11328
rect 5080 11144 5132 11150
rect 5078 11112 5080 11121
rect 5132 11112 5134 11121
rect 5078 11047 5134 11056
rect 4896 10804 4948 10810
rect 4896 10746 4948 10752
rect 4988 10804 5040 10810
rect 4988 10746 5040 10752
rect 4712 10736 4764 10742
rect 4712 10678 4764 10684
rect 4804 10736 4856 10742
rect 4804 10678 4856 10684
rect 4540 10526 4660 10554
rect 4540 7886 4568 10526
rect 4712 9920 4764 9926
rect 4632 9880 4712 9908
rect 4632 8974 4660 9880
rect 4712 9862 4764 9868
rect 4816 9738 4844 10678
rect 4908 9926 4936 10746
rect 5184 10690 5212 11698
rect 5000 10662 5212 10690
rect 5276 10690 5304 11834
rect 5368 11801 5396 12406
rect 5460 12238 5488 12786
rect 5644 12442 5672 12786
rect 5632 12436 5684 12442
rect 5632 12378 5684 12384
rect 5448 12232 5500 12238
rect 5448 12174 5500 12180
rect 5632 12164 5684 12170
rect 5632 12106 5684 12112
rect 5448 11892 5500 11898
rect 5448 11834 5500 11840
rect 5354 11792 5410 11801
rect 5354 11727 5410 11736
rect 5460 11676 5488 11834
rect 5368 11648 5488 11676
rect 5368 10810 5396 11648
rect 5540 11552 5592 11558
rect 5540 11494 5592 11500
rect 5448 11144 5500 11150
rect 5448 11086 5500 11092
rect 5460 10962 5488 11086
rect 5552 11064 5580 11494
rect 5644 11122 5672 12106
rect 5736 11558 5764 13670
rect 5828 13297 5856 13806
rect 5906 13767 5962 13776
rect 5814 13288 5870 13297
rect 5814 13223 5870 13232
rect 5828 12442 5856 13223
rect 5816 12436 5868 12442
rect 5816 12378 5868 12384
rect 5828 12345 5856 12378
rect 5814 12336 5870 12345
rect 5920 12306 5948 13767
rect 6012 12306 6040 14418
rect 6104 13569 6132 18702
rect 6196 17270 6224 19200
rect 8576 18284 8628 18290
rect 8576 18226 8628 18232
rect 6736 18216 6788 18222
rect 6366 18184 6422 18193
rect 6736 18158 6788 18164
rect 6366 18119 6422 18128
rect 6184 17264 6236 17270
rect 6184 17206 6236 17212
rect 6276 16992 6328 16998
rect 6276 16934 6328 16940
rect 6184 14612 6236 14618
rect 6184 14554 6236 14560
rect 6090 13560 6146 13569
rect 6090 13495 6146 13504
rect 6104 13394 6132 13495
rect 6092 13388 6144 13394
rect 6092 13330 6144 13336
rect 6196 13297 6224 14554
rect 6288 13734 6316 16934
rect 6380 13938 6408 18119
rect 6550 16552 6606 16561
rect 6550 16487 6606 16496
rect 6564 16114 6592 16487
rect 6552 16108 6604 16114
rect 6552 16050 6604 16056
rect 6644 16108 6696 16114
rect 6644 16050 6696 16056
rect 6460 16040 6512 16046
rect 6460 15982 6512 15988
rect 6472 15570 6500 15982
rect 6460 15564 6512 15570
rect 6460 15506 6512 15512
rect 6552 15428 6604 15434
rect 6552 15370 6604 15376
rect 6564 14550 6592 15370
rect 6656 15337 6684 16050
rect 6642 15328 6698 15337
rect 6642 15263 6698 15272
rect 6552 14544 6604 14550
rect 6552 14486 6604 14492
rect 6748 14056 6776 18158
rect 8208 17604 8260 17610
rect 8208 17546 8260 17552
rect 7610 17436 7918 17445
rect 7610 17434 7616 17436
rect 7672 17434 7696 17436
rect 7752 17434 7776 17436
rect 7832 17434 7856 17436
rect 7912 17434 7918 17436
rect 7672 17382 7674 17434
rect 7854 17382 7856 17434
rect 7610 17380 7616 17382
rect 7672 17380 7696 17382
rect 7752 17380 7776 17382
rect 7832 17380 7856 17382
rect 7912 17380 7918 17382
rect 7470 17368 7526 17377
rect 7610 17371 7918 17380
rect 7470 17303 7526 17312
rect 7380 17196 7432 17202
rect 7380 17138 7432 17144
rect 6950 16892 7258 16901
rect 6950 16890 6956 16892
rect 7012 16890 7036 16892
rect 7092 16890 7116 16892
rect 7172 16890 7196 16892
rect 7252 16890 7258 16892
rect 7012 16838 7014 16890
rect 7194 16838 7196 16890
rect 6950 16836 6956 16838
rect 7012 16836 7036 16838
rect 7092 16836 7116 16838
rect 7172 16836 7196 16838
rect 7252 16836 7258 16838
rect 6950 16827 7258 16836
rect 7392 16182 7420 17138
rect 7484 16833 7512 17303
rect 7470 16824 7526 16833
rect 7470 16759 7526 16768
rect 8116 16788 8168 16794
rect 8116 16730 8168 16736
rect 7610 16348 7918 16357
rect 7610 16346 7616 16348
rect 7672 16346 7696 16348
rect 7752 16346 7776 16348
rect 7832 16346 7856 16348
rect 7912 16346 7918 16348
rect 7672 16294 7674 16346
rect 7854 16294 7856 16346
rect 7610 16292 7616 16294
rect 7672 16292 7696 16294
rect 7752 16292 7776 16294
rect 7832 16292 7856 16294
rect 7912 16292 7918 16294
rect 7470 16280 7526 16289
rect 7610 16283 7918 16292
rect 7470 16215 7526 16224
rect 7380 16176 7432 16182
rect 7380 16118 7432 16124
rect 7012 16108 7064 16114
rect 7012 16050 7064 16056
rect 7024 16017 7052 16050
rect 7010 16008 7066 16017
rect 7010 15943 7066 15952
rect 7380 15904 7432 15910
rect 7378 15872 7380 15881
rect 7432 15872 7434 15881
rect 6950 15804 7258 15813
rect 7378 15807 7434 15816
rect 6950 15802 6956 15804
rect 7012 15802 7036 15804
rect 7092 15802 7116 15804
rect 7172 15802 7196 15804
rect 7252 15802 7258 15804
rect 7012 15750 7014 15802
rect 7194 15750 7196 15802
rect 6950 15748 6956 15750
rect 7012 15748 7036 15750
rect 7092 15748 7116 15750
rect 7172 15748 7196 15750
rect 7252 15748 7258 15750
rect 6950 15739 7258 15748
rect 7484 15745 7512 16215
rect 7840 16108 7892 16114
rect 7840 16050 7892 16056
rect 7748 16040 7800 16046
rect 7748 15982 7800 15988
rect 7470 15736 7526 15745
rect 7470 15671 7526 15680
rect 7288 15632 7340 15638
rect 6918 15600 6974 15609
rect 7288 15574 7340 15580
rect 6918 15535 6974 15544
rect 6932 15502 6960 15535
rect 6920 15496 6972 15502
rect 6920 15438 6972 15444
rect 6950 14716 7258 14725
rect 6950 14714 6956 14716
rect 7012 14714 7036 14716
rect 7092 14714 7116 14716
rect 7172 14714 7196 14716
rect 7252 14714 7258 14716
rect 7012 14662 7014 14714
rect 7194 14662 7196 14714
rect 6950 14660 6956 14662
rect 7012 14660 7036 14662
rect 7092 14660 7116 14662
rect 7172 14660 7196 14662
rect 7252 14660 7258 14662
rect 6950 14651 7258 14660
rect 6564 14028 6776 14056
rect 6368 13932 6420 13938
rect 6368 13874 6420 13880
rect 6460 13932 6512 13938
rect 6460 13874 6512 13880
rect 6472 13841 6500 13874
rect 6458 13832 6514 13841
rect 6458 13767 6514 13776
rect 6276 13728 6328 13734
rect 6276 13670 6328 13676
rect 6458 13560 6514 13569
rect 6458 13495 6514 13504
rect 6472 13394 6500 13495
rect 6460 13388 6512 13394
rect 6460 13330 6512 13336
rect 6276 13320 6328 13326
rect 6182 13288 6238 13297
rect 6092 13252 6144 13258
rect 6276 13262 6328 13268
rect 6182 13223 6238 13232
rect 6092 13194 6144 13200
rect 5814 12271 5870 12280
rect 5908 12300 5960 12306
rect 5908 12242 5960 12248
rect 6000 12300 6052 12306
rect 6000 12242 6052 12248
rect 6104 12050 6132 13194
rect 6182 12880 6238 12889
rect 6182 12815 6238 12824
rect 6196 12238 6224 12815
rect 6184 12232 6236 12238
rect 6184 12174 6236 12180
rect 5920 12022 6132 12050
rect 5920 11744 5948 12022
rect 5828 11716 5948 11744
rect 5998 11792 6054 11801
rect 5998 11727 6054 11736
rect 5724 11552 5776 11558
rect 5724 11494 5776 11500
rect 5722 11384 5778 11393
rect 5722 11319 5778 11328
rect 5736 11218 5764 11319
rect 5828 11257 5856 11716
rect 5906 11656 5962 11665
rect 5906 11591 5962 11600
rect 5814 11248 5870 11257
rect 5724 11212 5776 11218
rect 5814 11183 5870 11192
rect 5724 11154 5776 11160
rect 5920 11132 5948 11591
rect 6012 11354 6040 11727
rect 6092 11620 6144 11626
rect 6092 11562 6144 11568
rect 6000 11348 6052 11354
rect 6000 11290 6052 11296
rect 6000 11144 6052 11150
rect 5644 11094 5764 11122
rect 5920 11104 6000 11132
rect 5552 11036 5672 11064
rect 5460 10934 5580 10962
rect 5356 10804 5408 10810
rect 5356 10746 5408 10752
rect 5448 10804 5500 10810
rect 5448 10746 5500 10752
rect 5460 10713 5488 10746
rect 5446 10704 5502 10713
rect 5276 10662 5396 10690
rect 5000 10266 5028 10662
rect 5172 10600 5224 10606
rect 5092 10560 5172 10588
rect 4988 10260 5040 10266
rect 4988 10202 5040 10208
rect 4986 10160 5042 10169
rect 4986 10095 5042 10104
rect 5000 9994 5028 10095
rect 4988 9988 5040 9994
rect 4988 9930 5040 9936
rect 4896 9920 4948 9926
rect 4896 9862 4948 9868
rect 4816 9710 5028 9738
rect 4802 9616 4858 9625
rect 4802 9551 4858 9560
rect 4816 9330 4844 9551
rect 4894 9480 4950 9489
rect 4894 9415 4950 9424
rect 4724 9302 4844 9330
rect 4620 8968 4672 8974
rect 4620 8910 4672 8916
rect 4632 8265 4660 8910
rect 4724 8566 4752 9302
rect 4908 8922 4936 9415
rect 4816 8894 4936 8922
rect 4712 8560 4764 8566
rect 4712 8502 4764 8508
rect 4618 8256 4674 8265
rect 4618 8191 4674 8200
rect 4620 8084 4672 8090
rect 4620 8026 4672 8032
rect 4528 7880 4580 7886
rect 4528 7822 4580 7828
rect 4528 7336 4580 7342
rect 4528 7278 4580 7284
rect 4436 6792 4488 6798
rect 4436 6734 4488 6740
rect 4434 6624 4490 6633
rect 4434 6559 4490 6568
rect 4448 6390 4476 6559
rect 4436 6384 4488 6390
rect 4436 6326 4488 6332
rect 4436 6248 4488 6254
rect 4436 6190 4488 6196
rect 3976 5228 4028 5234
rect 3976 5170 4028 5176
rect 4160 5228 4212 5234
rect 4344 5228 4396 5234
rect 4160 5170 4212 5176
rect 4264 5188 4344 5216
rect 4068 5160 4120 5166
rect 4068 5102 4120 5108
rect 3974 4992 4030 5001
rect 3974 4927 4030 4936
rect 3988 4622 4016 4927
rect 3976 4616 4028 4622
rect 3976 4558 4028 4564
rect 3884 4276 3936 4282
rect 3884 4218 3936 4224
rect 3884 4140 3936 4146
rect 3884 4082 3936 4088
rect 3896 4049 3924 4082
rect 3882 4040 3938 4049
rect 3882 3975 3938 3984
rect 3884 2916 3936 2922
rect 3884 2858 3936 2864
rect 3424 2644 3476 2650
rect 3424 2586 3476 2592
rect 3792 2644 3844 2650
rect 3792 2586 3844 2592
rect 3332 2372 3384 2378
rect 3332 2314 3384 2320
rect 3238 2136 3294 2145
rect 3238 2071 3294 2080
rect 3148 944 3200 950
rect 3148 886 3200 892
rect 3344 800 3372 2314
rect 3330 0 3386 800
rect 3896 513 3924 2858
rect 3976 2848 4028 2854
rect 3976 2790 4028 2796
rect 3988 542 4016 2790
rect 4080 1970 4108 5102
rect 4160 5092 4212 5098
rect 4160 5034 4212 5040
rect 4172 4622 4200 5034
rect 4264 4758 4292 5188
rect 4344 5170 4396 5176
rect 4344 5024 4396 5030
rect 4344 4966 4396 4972
rect 4252 4752 4304 4758
rect 4252 4694 4304 4700
rect 4160 4616 4212 4622
rect 4160 4558 4212 4564
rect 4264 4146 4292 4694
rect 4356 4554 4384 4966
rect 4448 4690 4476 6190
rect 4540 5710 4568 7278
rect 4632 6202 4660 8026
rect 4724 7546 4752 8502
rect 4816 8362 4844 8894
rect 4896 8832 4948 8838
rect 4896 8774 4948 8780
rect 4804 8356 4856 8362
rect 4804 8298 4856 8304
rect 4712 7540 4764 7546
rect 4712 7482 4764 7488
rect 4710 7304 4766 7313
rect 4710 7239 4766 7248
rect 4724 6610 4752 7239
rect 4816 6730 4844 8298
rect 4908 8265 4936 8774
rect 4894 8256 4950 8265
rect 4894 8191 4950 8200
rect 4896 7472 4948 7478
rect 4896 7414 4948 7420
rect 4804 6724 4856 6730
rect 4804 6666 4856 6672
rect 4908 6633 4936 7414
rect 4894 6624 4950 6633
rect 4724 6582 4844 6610
rect 4632 6174 4752 6202
rect 4620 6112 4672 6118
rect 4620 6054 4672 6060
rect 4528 5704 4580 5710
rect 4528 5646 4580 5652
rect 4632 5556 4660 6054
rect 4540 5528 4660 5556
rect 4436 4684 4488 4690
rect 4436 4626 4488 4632
rect 4344 4548 4396 4554
rect 4344 4490 4396 4496
rect 4356 4146 4384 4490
rect 4448 4282 4476 4626
rect 4436 4276 4488 4282
rect 4436 4218 4488 4224
rect 4252 4140 4304 4146
rect 4252 4082 4304 4088
rect 4344 4140 4396 4146
rect 4344 4082 4396 4088
rect 4344 4004 4396 4010
rect 4344 3946 4396 3952
rect 4356 3913 4384 3946
rect 4342 3904 4398 3913
rect 4342 3839 4398 3848
rect 4356 3534 4384 3839
rect 4540 3652 4568 5528
rect 4724 5386 4752 6174
rect 4816 5778 4844 6582
rect 4894 6559 4950 6568
rect 4896 6384 4948 6390
rect 4896 6326 4948 6332
rect 4908 6225 4936 6326
rect 4894 6216 4950 6225
rect 4894 6151 4950 6160
rect 5000 6118 5028 9710
rect 5092 9178 5120 10560
rect 5172 10542 5224 10548
rect 5264 10600 5316 10606
rect 5264 10542 5316 10548
rect 5172 10056 5224 10062
rect 5172 9998 5224 10004
rect 5184 9518 5212 9998
rect 5276 9761 5304 10542
rect 5368 10198 5396 10662
rect 5446 10639 5502 10648
rect 5448 10600 5500 10606
rect 5448 10542 5500 10548
rect 5356 10192 5408 10198
rect 5356 10134 5408 10140
rect 5356 9988 5408 9994
rect 5356 9930 5408 9936
rect 5262 9752 5318 9761
rect 5262 9687 5318 9696
rect 5172 9512 5224 9518
rect 5170 9480 5172 9489
rect 5224 9480 5226 9489
rect 5170 9415 5226 9424
rect 5172 9376 5224 9382
rect 5172 9318 5224 9324
rect 5080 9172 5132 9178
rect 5080 9114 5132 9120
rect 5080 8968 5132 8974
rect 5080 8910 5132 8916
rect 5092 8401 5120 8910
rect 5078 8392 5134 8401
rect 5078 8327 5134 8336
rect 5080 8288 5132 8294
rect 5080 8230 5132 8236
rect 5092 6662 5120 8230
rect 5080 6656 5132 6662
rect 5080 6598 5132 6604
rect 5080 6316 5132 6322
rect 5080 6258 5132 6264
rect 4988 6112 5040 6118
rect 4988 6054 5040 6060
rect 4804 5772 4856 5778
rect 4804 5714 4856 5720
rect 4896 5772 4948 5778
rect 4896 5714 4948 5720
rect 4632 5358 4752 5386
rect 4632 4146 4660 5358
rect 4908 5284 4936 5714
rect 4724 5256 4936 5284
rect 4724 4690 4752 5256
rect 4988 5228 5040 5234
rect 4908 5188 4988 5216
rect 4804 5092 4856 5098
rect 4804 5034 4856 5040
rect 4816 4729 4844 5034
rect 4802 4720 4858 4729
rect 4712 4684 4764 4690
rect 4802 4655 4858 4664
rect 4712 4626 4764 4632
rect 4710 4584 4766 4593
rect 4710 4519 4712 4528
rect 4764 4519 4766 4528
rect 4712 4490 4764 4496
rect 4620 4140 4672 4146
rect 4620 4082 4672 4088
rect 4632 3777 4660 4082
rect 4804 4072 4856 4078
rect 4804 4014 4856 4020
rect 4618 3768 4674 3777
rect 4618 3703 4674 3712
rect 4540 3624 4660 3652
rect 4160 3528 4212 3534
rect 4160 3470 4212 3476
rect 4344 3528 4396 3534
rect 4528 3528 4580 3534
rect 4344 3470 4396 3476
rect 4526 3496 4528 3505
rect 4580 3496 4582 3505
rect 4068 1964 4120 1970
rect 4068 1906 4120 1912
rect 4172 1018 4200 3470
rect 4526 3431 4582 3440
rect 4252 2984 4304 2990
rect 4252 2926 4304 2932
rect 4264 2446 4292 2926
rect 4252 2440 4304 2446
rect 4252 2382 4304 2388
rect 4540 2310 4568 3431
rect 4528 2304 4580 2310
rect 4528 2246 4580 2252
rect 4632 1290 4660 3624
rect 4620 1284 4672 1290
rect 4620 1226 4672 1232
rect 4816 1193 4844 4014
rect 4908 3942 4936 5188
rect 4988 5170 5040 5176
rect 5092 4978 5120 6258
rect 5184 5234 5212 9318
rect 5368 9194 5396 9930
rect 5276 9166 5396 9194
rect 5276 8974 5304 9166
rect 5264 8968 5316 8974
rect 5356 8968 5408 8974
rect 5264 8910 5316 8916
rect 5354 8936 5356 8945
rect 5408 8936 5410 8945
rect 5354 8871 5410 8880
rect 5356 8832 5408 8838
rect 5262 8800 5318 8809
rect 5356 8774 5408 8780
rect 5262 8735 5318 8744
rect 5276 8634 5304 8735
rect 5264 8628 5316 8634
rect 5264 8570 5316 8576
rect 5262 8528 5318 8537
rect 5262 8463 5318 8472
rect 5276 8430 5304 8463
rect 5264 8424 5316 8430
rect 5264 8366 5316 8372
rect 5262 8120 5318 8129
rect 5262 8055 5264 8064
rect 5316 8055 5318 8064
rect 5264 8026 5316 8032
rect 5264 7540 5316 7546
rect 5264 7482 5316 7488
rect 5276 5574 5304 7482
rect 5264 5568 5316 5574
rect 5264 5510 5316 5516
rect 5172 5228 5224 5234
rect 5172 5170 5224 5176
rect 5170 5128 5226 5137
rect 5170 5063 5226 5072
rect 5264 5092 5316 5098
rect 5000 4950 5120 4978
rect 5000 4049 5028 4950
rect 5080 4820 5132 4826
rect 5080 4762 5132 4768
rect 5092 4604 5120 4762
rect 5184 4758 5212 5063
rect 5264 5034 5316 5040
rect 5172 4752 5224 4758
rect 5172 4694 5224 4700
rect 5276 4604 5304 5034
rect 5092 4576 5304 4604
rect 5080 4276 5132 4282
rect 5080 4218 5132 4224
rect 5172 4276 5224 4282
rect 5172 4218 5224 4224
rect 4986 4040 5042 4049
rect 4986 3975 5042 3984
rect 4896 3936 4948 3942
rect 4896 3878 4948 3884
rect 4986 3904 5042 3913
rect 4986 3839 5042 3848
rect 4896 3460 4948 3466
rect 4896 3402 4948 3408
rect 4908 2854 4936 3402
rect 5000 3097 5028 3839
rect 4986 3088 5042 3097
rect 4986 3023 5042 3032
rect 4896 2848 4948 2854
rect 4896 2790 4948 2796
rect 5000 2514 5028 3023
rect 5092 2922 5120 4218
rect 5184 3126 5212 4218
rect 5276 4146 5304 4576
rect 5264 4140 5316 4146
rect 5264 4082 5316 4088
rect 5264 3528 5316 3534
rect 5264 3470 5316 3476
rect 5172 3120 5224 3126
rect 5172 3062 5224 3068
rect 5080 2916 5132 2922
rect 5080 2858 5132 2864
rect 4988 2508 5040 2514
rect 4988 2450 5040 2456
rect 4802 1184 4858 1193
rect 4802 1119 4858 1128
rect 4160 1012 4212 1018
rect 4160 954 4212 960
rect 5184 814 5212 3062
rect 5172 808 5224 814
rect 5172 750 5224 756
rect 5276 678 5304 3470
rect 5368 2774 5396 8774
rect 5460 4826 5488 10542
rect 5552 8294 5580 10934
rect 5644 9994 5672 11036
rect 5736 10470 5764 11094
rect 6000 11086 6052 11092
rect 6000 10668 6052 10674
rect 5920 10628 6000 10656
rect 5920 10538 5948 10628
rect 6000 10610 6052 10616
rect 6104 10606 6132 11562
rect 6182 11520 6238 11529
rect 6182 11455 6238 11464
rect 6196 11150 6224 11455
rect 6184 11144 6236 11150
rect 6184 11086 6236 11092
rect 6182 10976 6238 10985
rect 6288 10962 6316 13262
rect 6366 13016 6422 13025
rect 6564 12968 6592 14028
rect 7300 13977 7328 15574
rect 7760 15502 7788 15982
rect 7748 15496 7800 15502
rect 7748 15438 7800 15444
rect 7852 15434 7880 16050
rect 8024 15904 8076 15910
rect 8024 15846 8076 15852
rect 8036 15502 8064 15846
rect 8024 15496 8076 15502
rect 8024 15438 8076 15444
rect 7840 15428 7892 15434
rect 7840 15370 7892 15376
rect 7472 15360 7524 15366
rect 7472 15302 7524 15308
rect 7286 13968 7342 13977
rect 6644 13932 6696 13938
rect 7286 13903 7342 13912
rect 6644 13874 6696 13880
rect 6366 12951 6422 12960
rect 6380 12617 6408 12951
rect 6472 12940 6592 12968
rect 6366 12608 6422 12617
rect 6366 12543 6422 12552
rect 6366 12200 6422 12209
rect 6366 12135 6422 12144
rect 6380 11830 6408 12135
rect 6368 11824 6420 11830
rect 6368 11766 6420 11772
rect 6472 11626 6500 12940
rect 6550 12880 6606 12889
rect 6550 12815 6552 12824
rect 6604 12815 6606 12824
rect 6552 12786 6604 12792
rect 6550 12744 6606 12753
rect 6550 12679 6606 12688
rect 6564 12170 6592 12679
rect 6552 12164 6604 12170
rect 6552 12106 6604 12112
rect 6460 11620 6512 11626
rect 6460 11562 6512 11568
rect 6552 11620 6604 11626
rect 6552 11562 6604 11568
rect 6368 11552 6420 11558
rect 6368 11494 6420 11500
rect 6380 11064 6408 11494
rect 6380 11036 6500 11064
rect 6472 10985 6500 11036
rect 6458 10976 6514 10985
rect 6288 10934 6408 10962
rect 6182 10911 6238 10920
rect 6092 10600 6144 10606
rect 5998 10568 6054 10577
rect 5908 10532 5960 10538
rect 6092 10542 6144 10548
rect 5998 10503 6000 10512
rect 5908 10474 5960 10480
rect 6052 10503 6054 10512
rect 6000 10474 6052 10480
rect 5724 10464 5776 10470
rect 5776 10424 5856 10452
rect 5724 10406 5776 10412
rect 5632 9988 5684 9994
rect 5632 9930 5684 9936
rect 5724 9920 5776 9926
rect 5724 9862 5776 9868
rect 5632 9580 5684 9586
rect 5632 9522 5684 9528
rect 5540 8288 5592 8294
rect 5540 8230 5592 8236
rect 5540 7268 5592 7274
rect 5540 7210 5592 7216
rect 5552 6458 5580 7210
rect 5540 6452 5592 6458
rect 5540 6394 5592 6400
rect 5540 6180 5592 6186
rect 5540 6122 5592 6128
rect 5448 4820 5500 4826
rect 5448 4762 5500 4768
rect 5552 4622 5580 6122
rect 5644 5234 5672 9522
rect 5736 8498 5764 9862
rect 5724 8492 5776 8498
rect 5724 8434 5776 8440
rect 5736 7002 5764 8434
rect 5724 6996 5776 7002
rect 5724 6938 5776 6944
rect 5828 6934 5856 10424
rect 6090 10024 6146 10033
rect 6090 9959 6146 9968
rect 5908 9716 5960 9722
rect 5908 9658 5960 9664
rect 5816 6928 5868 6934
rect 5722 6896 5778 6905
rect 5816 6870 5868 6876
rect 5722 6831 5778 6840
rect 5736 6322 5764 6831
rect 5816 6724 5868 6730
rect 5816 6666 5868 6672
rect 5724 6316 5776 6322
rect 5724 6258 5776 6264
rect 5828 5953 5856 6666
rect 5814 5944 5870 5953
rect 5814 5879 5870 5888
rect 5816 5568 5868 5574
rect 5816 5510 5868 5516
rect 5722 5264 5778 5273
rect 5632 5228 5684 5234
rect 5722 5199 5778 5208
rect 5632 5170 5684 5176
rect 5540 4616 5592 4622
rect 5446 4584 5502 4593
rect 5540 4558 5592 4564
rect 5446 4519 5502 4528
rect 5460 4185 5488 4519
rect 5446 4176 5502 4185
rect 5446 4111 5502 4120
rect 5460 4078 5488 4111
rect 5552 4078 5580 4558
rect 5448 4072 5500 4078
rect 5448 4014 5500 4020
rect 5540 4072 5592 4078
rect 5540 4014 5592 4020
rect 5448 3936 5500 3942
rect 5448 3878 5500 3884
rect 5460 3738 5488 3878
rect 5448 3732 5500 3738
rect 5448 3674 5500 3680
rect 5644 3670 5672 5170
rect 5736 5030 5764 5199
rect 5724 5024 5776 5030
rect 5724 4966 5776 4972
rect 5828 4826 5856 5510
rect 5920 5302 5948 9658
rect 5998 9208 6054 9217
rect 5998 9143 6054 9152
rect 6012 8634 6040 9143
rect 6000 8628 6052 8634
rect 6000 8570 6052 8576
rect 6000 8424 6052 8430
rect 5998 8392 6000 8401
rect 6052 8392 6054 8401
rect 5998 8327 6054 8336
rect 6000 7880 6052 7886
rect 6000 7822 6052 7828
rect 6012 5778 6040 7822
rect 6104 6866 6132 9959
rect 6196 9722 6224 10911
rect 6274 10840 6330 10849
rect 6274 10775 6330 10784
rect 6288 10674 6316 10775
rect 6276 10668 6328 10674
rect 6276 10610 6328 10616
rect 6380 10418 6408 10934
rect 6458 10911 6514 10920
rect 6458 10704 6514 10713
rect 6458 10639 6514 10648
rect 6472 10577 6500 10639
rect 6458 10568 6514 10577
rect 6458 10503 6514 10512
rect 6564 10470 6592 11562
rect 6288 10390 6408 10418
rect 6460 10464 6512 10470
rect 6460 10406 6512 10412
rect 6552 10464 6604 10470
rect 6552 10406 6604 10412
rect 6184 9716 6236 9722
rect 6184 9658 6236 9664
rect 6184 9580 6236 9586
rect 6184 9522 6236 9528
rect 6092 6860 6144 6866
rect 6092 6802 6144 6808
rect 6090 6760 6146 6769
rect 6090 6695 6146 6704
rect 6000 5772 6052 5778
rect 6000 5714 6052 5720
rect 5908 5296 5960 5302
rect 5908 5238 5960 5244
rect 6104 5148 6132 6695
rect 6196 6644 6224 9522
rect 6288 8022 6316 10390
rect 6368 10124 6420 10130
rect 6368 10066 6420 10072
rect 6380 9722 6408 10066
rect 6472 10033 6500 10406
rect 6458 10024 6514 10033
rect 6458 9959 6514 9968
rect 6458 9752 6514 9761
rect 6368 9716 6420 9722
rect 6458 9687 6514 9696
rect 6368 9658 6420 9664
rect 6368 9512 6420 9518
rect 6368 9454 6420 9460
rect 6380 9353 6408 9454
rect 6366 9344 6422 9353
rect 6366 9279 6422 9288
rect 6368 8968 6420 8974
rect 6368 8910 6420 8916
rect 6276 8016 6328 8022
rect 6276 7958 6328 7964
rect 6288 7478 6316 7958
rect 6276 7472 6328 7478
rect 6276 7414 6328 7420
rect 6276 7336 6328 7342
rect 6276 7278 6328 7284
rect 6288 6769 6316 7278
rect 6274 6760 6330 6769
rect 6274 6695 6330 6704
rect 6196 6616 6316 6644
rect 6184 6316 6236 6322
rect 6184 6258 6236 6264
rect 5920 5120 6132 5148
rect 5816 4820 5868 4826
rect 5816 4762 5868 4768
rect 5920 4706 5948 5120
rect 6000 5024 6052 5030
rect 6000 4966 6052 4972
rect 5736 4678 5948 4706
rect 5632 3664 5684 3670
rect 5446 3632 5502 3641
rect 5632 3606 5684 3612
rect 5446 3567 5502 3576
rect 5460 3126 5488 3567
rect 5630 3496 5686 3505
rect 5540 3460 5592 3466
rect 5630 3431 5686 3440
rect 5540 3402 5592 3408
rect 5552 3369 5580 3402
rect 5644 3398 5672 3431
rect 5632 3392 5684 3398
rect 5538 3360 5594 3369
rect 5632 3334 5684 3340
rect 5538 3295 5594 3304
rect 5448 3120 5500 3126
rect 5448 3062 5500 3068
rect 5736 3058 5764 4678
rect 5814 4448 5870 4457
rect 5814 4383 5870 4392
rect 5828 4214 5856 4383
rect 5816 4208 5868 4214
rect 5816 4150 5868 4156
rect 5908 3936 5960 3942
rect 5906 3904 5908 3913
rect 5960 3904 5962 3913
rect 5906 3839 5962 3848
rect 6012 3720 6040 4966
rect 6092 4480 6144 4486
rect 6092 4422 6144 4428
rect 6104 4321 6132 4422
rect 6090 4312 6146 4321
rect 6090 4247 6146 4256
rect 5920 3692 6040 3720
rect 5816 3596 5868 3602
rect 5816 3538 5868 3544
rect 5724 3052 5776 3058
rect 5724 2994 5776 3000
rect 5368 2746 5488 2774
rect 5460 2650 5488 2746
rect 5448 2644 5500 2650
rect 5448 2586 5500 2592
rect 5736 1494 5764 2994
rect 5724 1488 5776 1494
rect 5724 1430 5776 1436
rect 5828 1086 5856 3538
rect 5920 3448 5948 3692
rect 6092 3528 6144 3534
rect 6090 3496 6092 3505
rect 6144 3496 6146 3505
rect 5920 3420 6040 3448
rect 6090 3431 6146 3440
rect 5816 1080 5868 1086
rect 5816 1022 5868 1028
rect 6012 882 6040 3420
rect 6090 1864 6146 1873
rect 6090 1799 6146 1808
rect 6104 1358 6132 1799
rect 6196 1358 6224 6258
rect 6288 6225 6316 6616
rect 6274 6216 6330 6225
rect 6274 6151 6330 6160
rect 6276 6112 6328 6118
rect 6276 6054 6328 6060
rect 6288 1630 6316 6054
rect 6380 3738 6408 8910
rect 6472 8498 6500 9687
rect 6564 8498 6592 10406
rect 6460 8492 6512 8498
rect 6460 8434 6512 8440
rect 6552 8492 6604 8498
rect 6552 8434 6604 8440
rect 6472 7585 6500 8434
rect 6458 7576 6514 7585
rect 6458 7511 6514 7520
rect 6564 7256 6592 8434
rect 6656 8265 6684 13874
rect 6736 13796 6788 13802
rect 6736 13738 6788 13744
rect 6748 13462 6776 13738
rect 6828 13728 6880 13734
rect 6828 13670 6880 13676
rect 6736 13456 6788 13462
rect 6736 13398 6788 13404
rect 6736 12844 6788 12850
rect 6736 12786 6788 12792
rect 6748 12753 6776 12786
rect 6734 12744 6790 12753
rect 6734 12679 6790 12688
rect 6840 12646 6868 13670
rect 6950 13628 7258 13637
rect 6950 13626 6956 13628
rect 7012 13626 7036 13628
rect 7092 13626 7116 13628
rect 7172 13626 7196 13628
rect 7252 13626 7258 13628
rect 7012 13574 7014 13626
rect 7194 13574 7196 13626
rect 6950 13572 6956 13574
rect 7012 13572 7036 13574
rect 7092 13572 7116 13574
rect 7172 13572 7196 13574
rect 7252 13572 7258 13574
rect 6950 13563 7258 13572
rect 7300 13394 7328 13903
rect 6920 13388 6972 13394
rect 6920 13330 6972 13336
rect 7288 13388 7340 13394
rect 7288 13330 7340 13336
rect 6736 12640 6788 12646
rect 6736 12582 6788 12588
rect 6828 12640 6880 12646
rect 6932 12628 6960 13330
rect 7194 13288 7250 13297
rect 7194 13223 7250 13232
rect 7012 13184 7064 13190
rect 7012 13126 7064 13132
rect 7024 12850 7052 13126
rect 7012 12844 7064 12850
rect 7012 12786 7064 12792
rect 7012 12640 7064 12646
rect 6932 12600 7012 12628
rect 6828 12582 6880 12588
rect 7208 12628 7236 13223
rect 7378 13152 7434 13161
rect 7378 13087 7434 13096
rect 7286 13016 7342 13025
rect 7392 12986 7420 13087
rect 7286 12951 7342 12960
rect 7380 12980 7432 12986
rect 7300 12832 7328 12951
rect 7484 12968 7512 15302
rect 7610 15260 7918 15269
rect 7610 15258 7616 15260
rect 7672 15258 7696 15260
rect 7752 15258 7776 15260
rect 7832 15258 7856 15260
rect 7912 15258 7918 15260
rect 7672 15206 7674 15258
rect 7854 15206 7856 15258
rect 7610 15204 7616 15206
rect 7672 15204 7696 15206
rect 7752 15204 7776 15206
rect 7832 15204 7856 15206
rect 7912 15204 7918 15206
rect 7610 15195 7918 15204
rect 8024 15088 8076 15094
rect 8024 15030 8076 15036
rect 7610 14172 7918 14181
rect 7610 14170 7616 14172
rect 7672 14170 7696 14172
rect 7752 14170 7776 14172
rect 7832 14170 7856 14172
rect 7912 14170 7918 14172
rect 7672 14118 7674 14170
rect 7854 14118 7856 14170
rect 7610 14116 7616 14118
rect 7672 14116 7696 14118
rect 7752 14116 7776 14118
rect 7832 14116 7856 14118
rect 7912 14116 7918 14118
rect 7610 14107 7918 14116
rect 8036 14056 8064 15030
rect 7944 14028 8064 14056
rect 7748 13932 7800 13938
rect 7748 13874 7800 13880
rect 7564 13728 7616 13734
rect 7564 13670 7616 13676
rect 7576 13297 7604 13670
rect 7760 13297 7788 13874
rect 7944 13734 7972 14028
rect 8128 14006 8156 16730
rect 8220 16114 8248 17546
rect 8588 16658 8616 18226
rect 8680 17270 8708 19200
rect 10232 18624 10284 18630
rect 10232 18566 10284 18572
rect 10874 18592 10930 18601
rect 9680 18420 9732 18426
rect 9680 18362 9732 18368
rect 9036 18080 9088 18086
rect 9036 18022 9088 18028
rect 8668 17264 8720 17270
rect 8668 17206 8720 17212
rect 8666 17096 8722 17105
rect 8666 17031 8722 17040
rect 8576 16652 8628 16658
rect 8576 16594 8628 16600
rect 8208 16108 8260 16114
rect 8208 16050 8260 16056
rect 8484 15700 8536 15706
rect 8484 15642 8536 15648
rect 8300 15496 8352 15502
rect 8300 15438 8352 15444
rect 8208 15156 8260 15162
rect 8208 15098 8260 15104
rect 8220 14657 8248 15098
rect 8206 14648 8262 14657
rect 8206 14583 8262 14592
rect 8312 14385 8340 15438
rect 8392 15428 8444 15434
rect 8392 15370 8444 15376
rect 8404 15026 8432 15370
rect 8496 15201 8524 15642
rect 8576 15360 8628 15366
rect 8576 15302 8628 15308
rect 8482 15192 8538 15201
rect 8482 15127 8538 15136
rect 8392 15020 8444 15026
rect 8392 14962 8444 14968
rect 8404 14618 8432 14962
rect 8496 14958 8524 15127
rect 8588 14958 8616 15302
rect 8484 14952 8536 14958
rect 8484 14894 8536 14900
rect 8576 14952 8628 14958
rect 8576 14894 8628 14900
rect 8484 14816 8536 14822
rect 8484 14758 8536 14764
rect 8392 14612 8444 14618
rect 8392 14554 8444 14560
rect 8298 14376 8354 14385
rect 8298 14311 8354 14320
rect 8116 14000 8168 14006
rect 8312 13988 8340 14311
rect 8116 13942 8168 13948
rect 8220 13960 8340 13988
rect 8024 13932 8076 13938
rect 8024 13874 8076 13880
rect 7932 13728 7984 13734
rect 7932 13670 7984 13676
rect 7930 13560 7986 13569
rect 7930 13495 7986 13504
rect 7944 13326 7972 13495
rect 7932 13320 7984 13326
rect 7562 13288 7618 13297
rect 7562 13223 7618 13232
rect 7746 13288 7802 13297
rect 7932 13262 7984 13268
rect 7746 13223 7802 13232
rect 7610 13084 7918 13093
rect 7610 13082 7616 13084
rect 7672 13082 7696 13084
rect 7752 13082 7776 13084
rect 7832 13082 7856 13084
rect 7912 13082 7918 13084
rect 7672 13030 7674 13082
rect 7854 13030 7856 13082
rect 7610 13028 7616 13030
rect 7672 13028 7696 13030
rect 7752 13028 7776 13030
rect 7832 13028 7856 13030
rect 7912 13028 7918 13030
rect 7610 13019 7918 13028
rect 7656 12980 7708 12986
rect 7484 12940 7656 12968
rect 7380 12922 7432 12928
rect 7656 12922 7708 12928
rect 7564 12844 7616 12850
rect 7300 12804 7512 12832
rect 7208 12600 7420 12628
rect 7484 12617 7512 12804
rect 7748 12844 7800 12850
rect 7616 12804 7748 12832
rect 7564 12786 7616 12792
rect 7748 12786 7800 12792
rect 7564 12708 7616 12714
rect 7748 12708 7800 12714
rect 7616 12668 7748 12696
rect 7564 12650 7616 12656
rect 7748 12650 7800 12656
rect 7012 12582 7064 12588
rect 6748 11626 6776 12582
rect 6840 12424 6868 12582
rect 6950 12540 7258 12549
rect 6950 12538 6956 12540
rect 7012 12538 7036 12540
rect 7092 12538 7116 12540
rect 7172 12538 7196 12540
rect 7252 12538 7258 12540
rect 7012 12486 7014 12538
rect 7194 12486 7196 12538
rect 6950 12484 6956 12486
rect 7012 12484 7036 12486
rect 7092 12484 7116 12486
rect 7172 12484 7196 12486
rect 7252 12484 7258 12486
rect 6950 12475 7258 12484
rect 6840 12396 7328 12424
rect 7300 12306 7328 12396
rect 7012 12300 7064 12306
rect 7012 12242 7064 12248
rect 7288 12300 7340 12306
rect 7392 12288 7420 12600
rect 7470 12608 7526 12617
rect 7470 12543 7526 12552
rect 7656 12436 7708 12442
rect 7656 12378 7708 12384
rect 7668 12345 7696 12378
rect 7654 12336 7710 12345
rect 7392 12260 7512 12288
rect 7654 12271 7710 12280
rect 7288 12242 7340 12248
rect 7024 11762 7052 12242
rect 7102 12200 7158 12209
rect 7102 12135 7158 12144
rect 7380 12164 7432 12170
rect 7012 11756 7064 11762
rect 6840 11716 7012 11744
rect 6736 11620 6788 11626
rect 6736 11562 6788 11568
rect 6734 11520 6790 11529
rect 6734 11455 6790 11464
rect 6748 11354 6776 11455
rect 6736 11348 6788 11354
rect 6736 11290 6788 11296
rect 6840 11150 6868 11716
rect 7012 11698 7064 11704
rect 7116 11665 7144 12135
rect 7380 12106 7432 12112
rect 7392 11898 7420 12106
rect 7380 11892 7432 11898
rect 7380 11834 7432 11840
rect 7288 11824 7340 11830
rect 7288 11766 7340 11772
rect 7102 11656 7158 11665
rect 7300 11642 7328 11766
rect 7380 11756 7432 11762
rect 7484 11744 7512 12260
rect 8036 12220 8064 13874
rect 8220 13462 8248 13960
rect 8208 13456 8260 13462
rect 8208 13398 8260 13404
rect 8298 13424 8354 13433
rect 8116 13388 8168 13394
rect 8298 13359 8354 13368
rect 8116 13330 8168 13336
rect 8128 12374 8156 13330
rect 8312 13326 8340 13359
rect 8300 13320 8352 13326
rect 8300 13262 8352 13268
rect 8208 13252 8260 13258
rect 8208 13194 8260 13200
rect 8220 12442 8248 13194
rect 8404 12850 8432 14554
rect 8496 13870 8524 14758
rect 8576 14544 8628 14550
rect 8576 14486 8628 14492
rect 8588 13977 8616 14486
rect 8680 14074 8708 17031
rect 8760 16992 8812 16998
rect 8760 16934 8812 16940
rect 8772 14770 8800 16934
rect 8852 16652 8904 16658
rect 8852 16594 8904 16600
rect 8864 15502 8892 16594
rect 9048 15502 9076 18022
rect 9692 17898 9720 18362
rect 9600 17870 9720 17898
rect 9600 17814 9628 17870
rect 9588 17808 9640 17814
rect 9588 17750 9640 17756
rect 9864 17740 9916 17746
rect 9864 17682 9916 17688
rect 9876 17542 9904 17682
rect 9772 17536 9824 17542
rect 9772 17478 9824 17484
rect 9864 17536 9916 17542
rect 9864 17478 9916 17484
rect 9496 17332 9548 17338
rect 9496 17274 9548 17280
rect 9126 17232 9182 17241
rect 9126 17167 9182 17176
rect 9140 16697 9168 17167
rect 9126 16688 9182 16697
rect 9126 16623 9182 16632
rect 9128 16176 9180 16182
rect 9128 16118 9180 16124
rect 8852 15496 8904 15502
rect 9036 15496 9088 15502
rect 8852 15438 8904 15444
rect 8942 15464 8998 15473
rect 8864 15337 8892 15438
rect 9140 15473 9168 16118
rect 9220 16108 9272 16114
rect 9220 16050 9272 16056
rect 9036 15438 9088 15444
rect 9126 15464 9182 15473
rect 8942 15399 8998 15408
rect 9126 15399 9182 15408
rect 8850 15328 8906 15337
rect 8850 15263 8906 15272
rect 8772 14742 8892 14770
rect 8760 14544 8812 14550
rect 8760 14486 8812 14492
rect 8668 14068 8720 14074
rect 8668 14010 8720 14016
rect 8574 13968 8630 13977
rect 8574 13903 8630 13912
rect 8668 13932 8720 13938
rect 8668 13874 8720 13880
rect 8484 13864 8536 13870
rect 8484 13806 8536 13812
rect 8484 13728 8536 13734
rect 8484 13670 8536 13676
rect 8496 13161 8524 13670
rect 8574 13288 8630 13297
rect 8574 13223 8630 13232
rect 8482 13152 8538 13161
rect 8482 13087 8538 13096
rect 8392 12844 8444 12850
rect 8392 12786 8444 12792
rect 8300 12776 8352 12782
rect 8300 12718 8352 12724
rect 8208 12436 8260 12442
rect 8208 12378 8260 12384
rect 8116 12368 8168 12374
rect 8116 12310 8168 12316
rect 8036 12192 8248 12220
rect 7610 11996 7918 12005
rect 7610 11994 7616 11996
rect 7672 11994 7696 11996
rect 7752 11994 7776 11996
rect 7832 11994 7856 11996
rect 7912 11994 7918 11996
rect 7672 11942 7674 11994
rect 7854 11942 7856 11994
rect 7610 11940 7616 11942
rect 7672 11940 7696 11942
rect 7752 11940 7776 11942
rect 7832 11940 7856 11942
rect 7912 11940 7918 11942
rect 7610 11931 7918 11940
rect 8022 11928 8078 11937
rect 7564 11892 7616 11898
rect 8022 11863 8078 11872
rect 7564 11834 7616 11840
rect 7432 11716 7512 11744
rect 7380 11698 7432 11704
rect 7300 11614 7420 11642
rect 7102 11591 7158 11600
rect 7392 11529 7420 11614
rect 7378 11520 7434 11529
rect 6950 11452 7258 11461
rect 7378 11455 7434 11464
rect 6950 11450 6956 11452
rect 7012 11450 7036 11452
rect 7092 11450 7116 11452
rect 7172 11450 7196 11452
rect 7252 11450 7258 11452
rect 7012 11398 7014 11450
rect 7194 11398 7196 11450
rect 6950 11396 6956 11398
rect 7012 11396 7036 11398
rect 7092 11396 7116 11398
rect 7172 11396 7196 11398
rect 7252 11396 7258 11398
rect 6950 11387 7258 11396
rect 7104 11348 7156 11354
rect 7576 11336 7604 11834
rect 7748 11756 7800 11762
rect 7748 11698 7800 11704
rect 7104 11290 7156 11296
rect 7208 11308 7604 11336
rect 7116 11218 7144 11290
rect 6920 11212 6972 11218
rect 6920 11154 6972 11160
rect 7104 11212 7156 11218
rect 7104 11154 7156 11160
rect 6828 11144 6880 11150
rect 6828 11086 6880 11092
rect 6736 11008 6788 11014
rect 6736 10950 6788 10956
rect 6748 8498 6776 10950
rect 6840 10849 6868 11086
rect 6932 10985 6960 11154
rect 7012 11076 7064 11082
rect 7012 11018 7064 11024
rect 6918 10976 6974 10985
rect 6918 10911 6974 10920
rect 6826 10840 6882 10849
rect 7024 10792 7052 11018
rect 6826 10775 6882 10784
rect 6932 10764 7052 10792
rect 6828 10668 6880 10674
rect 6932 10656 6960 10764
rect 6880 10628 6960 10656
rect 7010 10704 7066 10713
rect 7066 10662 7139 10690
rect 7208 10674 7236 11308
rect 7472 11212 7524 11218
rect 7472 11154 7524 11160
rect 7286 10976 7342 10985
rect 7286 10911 7342 10920
rect 7300 10674 7328 10911
rect 7484 10792 7512 11154
rect 7760 11082 7788 11698
rect 8036 11694 8064 11863
rect 7840 11688 7892 11694
rect 7840 11630 7892 11636
rect 8024 11688 8076 11694
rect 8024 11630 8076 11636
rect 7852 11082 7880 11630
rect 7932 11552 7984 11558
rect 7932 11494 7984 11500
rect 7944 11393 7972 11494
rect 7930 11384 7986 11393
rect 7930 11319 7986 11328
rect 8116 11280 8168 11286
rect 7930 11248 7986 11257
rect 8116 11222 8168 11228
rect 7930 11183 7986 11192
rect 7748 11076 7800 11082
rect 7748 11018 7800 11024
rect 7840 11076 7892 11082
rect 7840 11018 7892 11024
rect 7944 10996 7972 11183
rect 7944 10968 8064 10996
rect 7610 10908 7918 10917
rect 7610 10906 7616 10908
rect 7672 10906 7696 10908
rect 7752 10906 7776 10908
rect 7832 10906 7856 10908
rect 7912 10906 7918 10908
rect 7672 10854 7674 10906
rect 7854 10854 7856 10906
rect 7610 10852 7616 10854
rect 7672 10852 7696 10854
rect 7752 10852 7776 10854
rect 7832 10852 7856 10854
rect 7912 10852 7918 10854
rect 7610 10843 7918 10852
rect 7484 10764 7604 10792
rect 7470 10704 7526 10713
rect 7010 10639 7066 10648
rect 7111 10656 7139 10662
rect 7196 10668 7248 10674
rect 7111 10628 7144 10656
rect 6828 10610 6880 10616
rect 6840 9926 6868 10610
rect 7116 10538 7144 10628
rect 7196 10610 7248 10616
rect 7288 10668 7340 10674
rect 7470 10639 7526 10648
rect 7288 10610 7340 10616
rect 7104 10532 7156 10538
rect 7104 10474 7156 10480
rect 6950 10364 7258 10373
rect 6950 10362 6956 10364
rect 7012 10362 7036 10364
rect 7092 10362 7116 10364
rect 7172 10362 7196 10364
rect 7252 10362 7258 10364
rect 7012 10310 7014 10362
rect 7194 10310 7196 10362
rect 6950 10308 6956 10310
rect 7012 10308 7036 10310
rect 7092 10308 7116 10310
rect 7172 10308 7196 10310
rect 7252 10308 7258 10310
rect 6950 10299 7258 10308
rect 7300 10248 7328 10610
rect 7484 10606 7512 10639
rect 7472 10600 7524 10606
rect 7472 10542 7524 10548
rect 7470 10432 7526 10441
rect 7470 10367 7526 10376
rect 6932 10220 7328 10248
rect 6828 9920 6880 9926
rect 6828 9862 6880 9868
rect 6828 9648 6880 9654
rect 6828 9590 6880 9596
rect 6840 9382 6868 9590
rect 6932 9466 6960 10220
rect 7484 10180 7512 10367
rect 7392 10152 7512 10180
rect 7012 10124 7064 10130
rect 7392 10112 7420 10152
rect 7064 10084 7420 10112
rect 7012 10066 7064 10072
rect 7104 9988 7156 9994
rect 7104 9930 7156 9936
rect 7380 9988 7432 9994
rect 7576 9976 7604 10764
rect 7840 10736 7892 10742
rect 8036 10724 8064 10968
rect 7892 10696 8064 10724
rect 7840 10678 7892 10684
rect 7656 10668 7708 10674
rect 7656 10610 7708 10616
rect 7668 10470 7696 10610
rect 7748 10600 7800 10606
rect 7748 10542 7800 10548
rect 7656 10464 7708 10470
rect 7656 10406 7708 10412
rect 7654 10296 7710 10305
rect 7654 10231 7710 10240
rect 7380 9930 7432 9936
rect 7484 9948 7604 9976
rect 7116 9586 7144 9930
rect 7104 9580 7156 9586
rect 7104 9522 7156 9528
rect 6932 9438 7328 9466
rect 6828 9376 6880 9382
rect 6828 9318 6880 9324
rect 6950 9276 7258 9285
rect 6950 9274 6956 9276
rect 7012 9274 7036 9276
rect 7092 9274 7116 9276
rect 7172 9274 7196 9276
rect 7252 9274 7258 9276
rect 7012 9222 7014 9274
rect 7194 9222 7196 9274
rect 6950 9220 6956 9222
rect 7012 9220 7036 9222
rect 7092 9220 7116 9222
rect 7172 9220 7196 9222
rect 7252 9220 7258 9222
rect 6950 9211 7258 9220
rect 6828 9172 6880 9178
rect 6828 9114 6880 9120
rect 6840 8498 6868 9114
rect 7104 9036 7156 9042
rect 7104 8978 7156 8984
rect 7010 8664 7066 8673
rect 7116 8634 7144 8978
rect 7196 8832 7248 8838
rect 7196 8774 7248 8780
rect 7010 8599 7066 8608
rect 7104 8628 7156 8634
rect 6736 8492 6788 8498
rect 6736 8434 6788 8440
rect 6828 8492 6880 8498
rect 6828 8434 6880 8440
rect 6642 8256 6698 8265
rect 6642 8191 6698 8200
rect 6734 8120 6790 8129
rect 6734 8055 6790 8064
rect 6840 8072 6868 8434
rect 7024 8294 7052 8599
rect 7104 8570 7156 8576
rect 7208 8412 7236 8774
rect 7300 8537 7328 9438
rect 7392 9353 7420 9930
rect 7378 9344 7434 9353
rect 7378 9279 7434 9288
rect 7378 9208 7434 9217
rect 7378 9143 7434 9152
rect 7392 9042 7420 9143
rect 7380 9036 7432 9042
rect 7380 8978 7432 8984
rect 7392 8945 7420 8978
rect 7378 8936 7434 8945
rect 7378 8871 7434 8880
rect 7378 8800 7434 8809
rect 7378 8735 7434 8744
rect 7286 8528 7342 8537
rect 7286 8463 7342 8472
rect 7208 8384 7328 8412
rect 7012 8288 7064 8294
rect 7012 8230 7064 8236
rect 6950 8188 7258 8197
rect 6950 8186 6956 8188
rect 7012 8186 7036 8188
rect 7092 8186 7116 8188
rect 7172 8186 7196 8188
rect 7252 8186 7258 8188
rect 7012 8134 7014 8186
rect 7194 8134 7196 8186
rect 6950 8132 6956 8134
rect 7012 8132 7036 8134
rect 7092 8132 7116 8134
rect 7172 8132 7196 8134
rect 7252 8132 7258 8134
rect 6950 8123 7258 8132
rect 7300 8072 7328 8384
rect 6748 7970 6776 8055
rect 6840 8044 6960 8072
rect 6644 7948 6696 7954
rect 6748 7942 6868 7970
rect 6644 7890 6696 7896
rect 6472 7228 6592 7256
rect 6472 6934 6500 7228
rect 6656 7154 6684 7890
rect 6736 7880 6788 7886
rect 6736 7822 6788 7828
rect 6564 7126 6684 7154
rect 6460 6928 6512 6934
rect 6460 6870 6512 6876
rect 6458 5808 6514 5817
rect 6458 5743 6514 5752
rect 6472 5710 6500 5743
rect 6460 5704 6512 5710
rect 6460 5646 6512 5652
rect 6460 5228 6512 5234
rect 6460 5170 6512 5176
rect 6472 4214 6500 5170
rect 6460 4208 6512 4214
rect 6460 4150 6512 4156
rect 6460 3936 6512 3942
rect 6460 3878 6512 3884
rect 6472 3777 6500 3878
rect 6458 3768 6514 3777
rect 6368 3732 6420 3738
rect 6458 3703 6514 3712
rect 6368 3674 6420 3680
rect 6564 3602 6592 7126
rect 6644 6792 6696 6798
rect 6642 6760 6644 6769
rect 6696 6760 6698 6769
rect 6642 6695 6698 6704
rect 6656 6322 6684 6695
rect 6644 6316 6696 6322
rect 6644 6258 6696 6264
rect 6642 6216 6698 6225
rect 6642 6151 6698 6160
rect 6656 5778 6684 6151
rect 6644 5772 6696 5778
rect 6644 5714 6696 5720
rect 6748 5658 6776 7822
rect 6840 5896 6868 7942
rect 6932 7342 6960 8044
rect 7208 8044 7328 8072
rect 7102 7984 7158 7993
rect 7208 7954 7236 8044
rect 7102 7919 7158 7928
rect 7196 7948 7248 7954
rect 7012 7744 7064 7750
rect 7012 7686 7064 7692
rect 6920 7336 6972 7342
rect 6920 7278 6972 7284
rect 7024 7274 7052 7686
rect 7116 7342 7144 7919
rect 7196 7890 7248 7896
rect 7288 7948 7340 7954
rect 7288 7890 7340 7896
rect 7196 7812 7248 7818
rect 7196 7754 7248 7760
rect 7208 7721 7236 7754
rect 7194 7712 7250 7721
rect 7194 7647 7250 7656
rect 7104 7336 7156 7342
rect 7104 7278 7156 7284
rect 7012 7268 7064 7274
rect 7012 7210 7064 7216
rect 6950 7100 7258 7109
rect 6950 7098 6956 7100
rect 7012 7098 7036 7100
rect 7092 7098 7116 7100
rect 7172 7098 7196 7100
rect 7252 7098 7258 7100
rect 7012 7046 7014 7098
rect 7194 7046 7196 7098
rect 6950 7044 6956 7046
rect 7012 7044 7036 7046
rect 7092 7044 7116 7046
rect 7172 7044 7196 7046
rect 7252 7044 7258 7046
rect 6950 7035 7258 7044
rect 7300 6984 7328 7890
rect 7116 6956 7328 6984
rect 7116 6254 7144 6956
rect 7392 6712 7420 8735
rect 7300 6684 7420 6712
rect 7196 6656 7248 6662
rect 7196 6598 7248 6604
rect 7208 6304 7236 6598
rect 7300 6497 7328 6684
rect 7378 6624 7434 6633
rect 7378 6559 7434 6568
rect 7286 6488 7342 6497
rect 7286 6423 7342 6432
rect 7288 6316 7340 6322
rect 7208 6276 7288 6304
rect 7288 6258 7340 6264
rect 7104 6248 7156 6254
rect 7104 6190 7156 6196
rect 6950 6012 7258 6021
rect 6950 6010 6956 6012
rect 7012 6010 7036 6012
rect 7092 6010 7116 6012
rect 7172 6010 7196 6012
rect 7252 6010 7258 6012
rect 7012 5958 7014 6010
rect 7194 5958 7196 6010
rect 6950 5956 6956 5958
rect 7012 5956 7036 5958
rect 7092 5956 7116 5958
rect 7172 5956 7196 5958
rect 7252 5956 7258 5958
rect 6950 5947 7258 5956
rect 7300 5896 7328 6258
rect 6840 5868 7144 5896
rect 7010 5808 7066 5817
rect 6828 5772 6880 5778
rect 7010 5743 7066 5752
rect 6828 5714 6880 5720
rect 6656 5630 6776 5658
rect 6656 4729 6684 5630
rect 6736 5568 6788 5574
rect 6734 5536 6736 5545
rect 6788 5536 6790 5545
rect 6734 5471 6790 5480
rect 6736 5024 6788 5030
rect 6734 4992 6736 5001
rect 6788 4992 6790 5001
rect 6734 4927 6790 4936
rect 6736 4820 6788 4826
rect 6736 4762 6788 4768
rect 6642 4720 6698 4729
rect 6642 4655 6698 4664
rect 6642 4448 6698 4457
rect 6642 4383 6698 4392
rect 6552 3596 6604 3602
rect 6552 3538 6604 3544
rect 6368 3460 6420 3466
rect 6368 3402 6420 3408
rect 6276 1624 6328 1630
rect 6276 1566 6328 1572
rect 6092 1352 6144 1358
rect 6092 1294 6144 1300
rect 6184 1352 6236 1358
rect 6184 1294 6236 1300
rect 6380 1154 6408 3402
rect 6656 3058 6684 4383
rect 6748 3194 6776 4762
rect 6840 4554 6868 5714
rect 7024 5166 7052 5743
rect 7116 5681 7144 5868
rect 7208 5868 7328 5896
rect 7102 5672 7158 5681
rect 7102 5607 7158 5616
rect 7012 5160 7064 5166
rect 7012 5102 7064 5108
rect 7208 5114 7236 5868
rect 7286 5536 7342 5545
rect 7286 5471 7342 5480
rect 7300 5370 7328 5471
rect 7288 5364 7340 5370
rect 7288 5306 7340 5312
rect 7300 5234 7328 5306
rect 7288 5228 7340 5234
rect 7288 5170 7340 5176
rect 7208 5086 7328 5114
rect 6950 4924 7258 4933
rect 6950 4922 6956 4924
rect 7012 4922 7036 4924
rect 7092 4922 7116 4924
rect 7172 4922 7196 4924
rect 7252 4922 7258 4924
rect 7012 4870 7014 4922
rect 7194 4870 7196 4922
rect 6950 4868 6956 4870
rect 7012 4868 7036 4870
rect 7092 4868 7116 4870
rect 7172 4868 7196 4870
rect 7252 4868 7258 4870
rect 6950 4859 7258 4868
rect 7012 4752 7064 4758
rect 7196 4752 7248 4758
rect 7064 4712 7196 4740
rect 7012 4694 7064 4700
rect 7196 4694 7248 4700
rect 7196 4616 7248 4622
rect 7196 4558 7248 4564
rect 6828 4548 6880 4554
rect 6828 4490 6880 4496
rect 7208 4185 7236 4558
rect 7194 4176 7250 4185
rect 7194 4111 7250 4120
rect 6950 3836 7258 3845
rect 6950 3834 6956 3836
rect 7012 3834 7036 3836
rect 7092 3834 7116 3836
rect 7172 3834 7196 3836
rect 7252 3834 7258 3836
rect 7012 3782 7014 3834
rect 7194 3782 7196 3834
rect 6950 3780 6956 3782
rect 7012 3780 7036 3782
rect 7092 3780 7116 3782
rect 7172 3780 7196 3782
rect 7252 3780 7258 3782
rect 6950 3771 7258 3780
rect 6932 3692 7236 3720
rect 6932 3534 6960 3692
rect 7208 3641 7236 3692
rect 7010 3632 7066 3641
rect 7010 3567 7066 3576
rect 7194 3632 7250 3641
rect 7300 3602 7328 5086
rect 7392 4826 7420 6559
rect 7484 5710 7512 9948
rect 7668 9926 7696 10231
rect 7760 10198 7788 10542
rect 8024 10464 8076 10470
rect 8024 10406 8076 10412
rect 7748 10192 7800 10198
rect 7748 10134 7800 10140
rect 7644 9920 7696 9926
rect 7644 9862 7696 9868
rect 7610 9820 7918 9829
rect 7610 9818 7616 9820
rect 7672 9818 7696 9820
rect 7752 9818 7776 9820
rect 7832 9818 7856 9820
rect 7912 9818 7918 9820
rect 7672 9766 7674 9818
rect 7854 9766 7856 9818
rect 7610 9764 7616 9766
rect 7672 9764 7696 9766
rect 7752 9764 7776 9766
rect 7832 9764 7856 9766
rect 7912 9764 7918 9766
rect 7610 9755 7918 9764
rect 8036 9704 8064 10406
rect 7852 9676 8064 9704
rect 7748 9580 7800 9586
rect 7748 9522 7800 9528
rect 7656 9512 7708 9518
rect 7656 9454 7708 9460
rect 7668 8945 7696 9454
rect 7760 9178 7788 9522
rect 7748 9172 7800 9178
rect 7748 9114 7800 9120
rect 7654 8936 7710 8945
rect 7654 8871 7710 8880
rect 7852 8838 7880 9676
rect 7932 9512 7984 9518
rect 7932 9454 7984 9460
rect 7944 8906 7972 9454
rect 8128 9160 8156 11222
rect 8220 10996 8248 12192
rect 8312 11064 8340 12718
rect 8392 12640 8444 12646
rect 8392 12582 8444 12588
rect 8404 11762 8432 12582
rect 8588 12288 8616 13223
rect 8496 12260 8616 12288
rect 8392 11756 8444 11762
rect 8392 11698 8444 11704
rect 8392 11620 8444 11626
rect 8496 11608 8524 12260
rect 8680 12220 8708 13874
rect 8444 11580 8524 11608
rect 8392 11562 8444 11568
rect 8312 11036 8432 11064
rect 8220 10968 8340 10996
rect 8208 10804 8260 10810
rect 8208 10746 8260 10752
rect 8220 10674 8248 10746
rect 8208 10668 8260 10674
rect 8208 10610 8260 10616
rect 8312 10470 8340 10968
rect 8300 10464 8352 10470
rect 8300 10406 8352 10412
rect 8206 10296 8262 10305
rect 8206 10231 8208 10240
rect 8260 10231 8262 10240
rect 8208 10202 8260 10208
rect 8206 9888 8262 9897
rect 8206 9823 8262 9832
rect 8220 9382 8248 9823
rect 8208 9376 8260 9382
rect 8404 9330 8432 11036
rect 8496 10962 8524 11580
rect 8588 12192 8708 12220
rect 8588 11558 8616 12192
rect 8772 12170 8800 14486
rect 8760 12164 8812 12170
rect 8680 12124 8760 12152
rect 8576 11552 8628 11558
rect 8576 11494 8628 11500
rect 8588 11218 8616 11494
rect 8576 11212 8628 11218
rect 8576 11154 8628 11160
rect 8496 10934 8632 10962
rect 8604 10724 8632 10934
rect 8588 10696 8632 10724
rect 8588 10690 8616 10696
rect 8208 9318 8260 9324
rect 8036 9132 8156 9160
rect 8312 9302 8432 9330
rect 8496 10662 8616 10690
rect 7932 8900 7984 8906
rect 7932 8842 7984 8848
rect 7840 8832 7892 8838
rect 7840 8774 7892 8780
rect 7610 8732 7918 8741
rect 7610 8730 7616 8732
rect 7672 8730 7696 8732
rect 7752 8730 7776 8732
rect 7832 8730 7856 8732
rect 7912 8730 7918 8732
rect 7672 8678 7674 8730
rect 7854 8678 7856 8730
rect 7610 8676 7616 8678
rect 7672 8676 7696 8678
rect 7752 8676 7776 8678
rect 7832 8676 7856 8678
rect 7912 8676 7918 8678
rect 7610 8667 7918 8676
rect 7656 8628 7708 8634
rect 7656 8570 7708 8576
rect 7748 8628 7800 8634
rect 7748 8570 7800 8576
rect 7668 8498 7696 8570
rect 7564 8492 7616 8498
rect 7564 8434 7616 8440
rect 7656 8492 7708 8498
rect 7656 8434 7708 8440
rect 7576 8265 7604 8434
rect 7562 8256 7618 8265
rect 7562 8191 7618 8200
rect 7562 8120 7618 8129
rect 7562 8055 7618 8064
rect 7576 7886 7604 8055
rect 7760 7993 7788 8570
rect 7840 8424 7892 8430
rect 7840 8366 7892 8372
rect 7746 7984 7802 7993
rect 7746 7919 7802 7928
rect 7852 7886 7880 8366
rect 7930 8256 7986 8265
rect 7930 8191 7986 8200
rect 7944 7954 7972 8191
rect 7932 7948 7984 7954
rect 7932 7890 7984 7896
rect 7564 7880 7616 7886
rect 7564 7822 7616 7828
rect 7840 7880 7892 7886
rect 7840 7822 7892 7828
rect 7610 7644 7918 7653
rect 7610 7642 7616 7644
rect 7672 7642 7696 7644
rect 7752 7642 7776 7644
rect 7832 7642 7856 7644
rect 7912 7642 7918 7644
rect 7672 7590 7674 7642
rect 7854 7590 7856 7642
rect 7610 7588 7616 7590
rect 7672 7588 7696 7590
rect 7752 7588 7776 7590
rect 7832 7588 7856 7590
rect 7912 7588 7918 7590
rect 7610 7579 7918 7588
rect 7564 7404 7616 7410
rect 7564 7346 7616 7352
rect 7576 7313 7604 7346
rect 7656 7336 7708 7342
rect 7562 7304 7618 7313
rect 7656 7278 7708 7284
rect 7562 7239 7618 7248
rect 7668 6798 7696 7278
rect 8036 7002 8064 9132
rect 8114 9072 8170 9081
rect 8114 9007 8116 9016
rect 8168 9007 8170 9016
rect 8116 8978 8168 8984
rect 8116 8900 8168 8906
rect 8116 8842 8168 8848
rect 8128 8294 8156 8842
rect 8208 8832 8260 8838
rect 8312 8809 8340 9302
rect 8392 9172 8444 9178
rect 8392 9114 8444 9120
rect 8208 8774 8260 8780
rect 8298 8800 8354 8809
rect 8116 8288 8168 8294
rect 8116 8230 8168 8236
rect 8128 7993 8156 8230
rect 8114 7984 8170 7993
rect 8114 7919 8170 7928
rect 8220 7886 8248 8774
rect 8298 8735 8354 8744
rect 8404 8673 8432 9114
rect 8390 8664 8446 8673
rect 8390 8599 8446 8608
rect 8298 7984 8354 7993
rect 8298 7919 8354 7928
rect 8208 7880 8260 7886
rect 8208 7822 8260 7828
rect 8116 7744 8168 7750
rect 8116 7686 8168 7692
rect 8128 7410 8156 7686
rect 8116 7404 8168 7410
rect 8116 7346 8168 7352
rect 8024 6996 8076 7002
rect 7944 6956 8024 6984
rect 7564 6792 7616 6798
rect 7562 6760 7564 6769
rect 7656 6792 7708 6798
rect 7616 6760 7618 6769
rect 7656 6734 7708 6740
rect 7562 6695 7618 6704
rect 7944 6662 7972 6956
rect 8024 6938 8076 6944
rect 8116 6996 8168 7002
rect 8116 6938 8168 6944
rect 8128 6798 8156 6938
rect 8220 6798 8248 7822
rect 8312 7478 8340 7919
rect 8392 7880 8444 7886
rect 8392 7822 8444 7828
rect 8404 7546 8432 7822
rect 8392 7540 8444 7546
rect 8392 7482 8444 7488
rect 8300 7472 8352 7478
rect 8300 7414 8352 7420
rect 8312 7177 8340 7414
rect 8392 7200 8444 7206
rect 8298 7168 8354 7177
rect 8392 7142 8444 7148
rect 8298 7103 8354 7112
rect 8404 6934 8432 7142
rect 8300 6928 8352 6934
rect 8300 6870 8352 6876
rect 8392 6928 8444 6934
rect 8392 6870 8444 6876
rect 8024 6792 8076 6798
rect 8024 6734 8076 6740
rect 8116 6792 8168 6798
rect 8116 6734 8168 6740
rect 8208 6792 8260 6798
rect 8312 6780 8340 6870
rect 8392 6792 8444 6798
rect 8312 6752 8392 6780
rect 8208 6734 8260 6740
rect 8392 6734 8444 6740
rect 7932 6656 7984 6662
rect 7932 6598 7984 6604
rect 7610 6556 7918 6565
rect 7610 6554 7616 6556
rect 7672 6554 7696 6556
rect 7752 6554 7776 6556
rect 7832 6554 7856 6556
rect 7912 6554 7918 6556
rect 7672 6502 7674 6554
rect 7854 6502 7856 6554
rect 7610 6500 7616 6502
rect 7672 6500 7696 6502
rect 7752 6500 7776 6502
rect 7832 6500 7856 6502
rect 7912 6500 7918 6502
rect 7610 6491 7918 6500
rect 7564 6452 7616 6458
rect 7564 6394 7616 6400
rect 7932 6452 7984 6458
rect 7932 6394 7984 6400
rect 7576 6254 7604 6394
rect 7656 6384 7708 6390
rect 7656 6326 7708 6332
rect 7564 6248 7616 6254
rect 7564 6190 7616 6196
rect 7668 6118 7696 6326
rect 7656 6112 7708 6118
rect 7656 6054 7708 6060
rect 7654 5944 7710 5953
rect 7654 5879 7710 5888
rect 7840 5908 7892 5914
rect 7668 5710 7696 5879
rect 7840 5850 7892 5856
rect 7472 5704 7524 5710
rect 7472 5646 7524 5652
rect 7656 5704 7708 5710
rect 7656 5646 7708 5652
rect 7852 5574 7880 5850
rect 7944 5574 7972 6394
rect 8036 6304 8064 6734
rect 8128 6458 8156 6734
rect 8208 6656 8260 6662
rect 8208 6598 8260 6604
rect 8300 6656 8352 6662
rect 8300 6598 8352 6604
rect 8116 6452 8168 6458
rect 8116 6394 8168 6400
rect 8220 6322 8248 6598
rect 8116 6316 8168 6322
rect 8036 6276 8116 6304
rect 8116 6258 8168 6264
rect 8208 6316 8260 6322
rect 8208 6258 8260 6264
rect 8116 6180 8168 6186
rect 8116 6122 8168 6128
rect 8022 6080 8078 6089
rect 8022 6015 8078 6024
rect 7840 5568 7892 5574
rect 7840 5510 7892 5516
rect 7932 5568 7984 5574
rect 7932 5510 7984 5516
rect 7610 5468 7918 5477
rect 7610 5466 7616 5468
rect 7672 5466 7696 5468
rect 7752 5466 7776 5468
rect 7832 5466 7856 5468
rect 7912 5466 7918 5468
rect 7672 5414 7674 5466
rect 7854 5414 7856 5466
rect 7610 5412 7616 5414
rect 7672 5412 7696 5414
rect 7752 5412 7776 5414
rect 7832 5412 7856 5414
rect 7912 5412 7918 5414
rect 7470 5400 7526 5409
rect 7610 5403 7918 5412
rect 7470 5335 7472 5344
rect 7524 5335 7526 5344
rect 7748 5364 7800 5370
rect 7472 5306 7524 5312
rect 7748 5306 7800 5312
rect 7472 5160 7524 5166
rect 7472 5102 7524 5108
rect 7380 4820 7432 4826
rect 7380 4762 7432 4768
rect 7378 4312 7434 4321
rect 7378 4247 7434 4256
rect 7194 3567 7250 3576
rect 7288 3596 7340 3602
rect 7024 3534 7052 3567
rect 7288 3538 7340 3544
rect 7392 3534 7420 4247
rect 7484 4146 7512 5102
rect 7760 4622 7788 5306
rect 7932 5228 7984 5234
rect 7932 5170 7984 5176
rect 7748 4616 7800 4622
rect 7944 4593 7972 5170
rect 8036 4622 8064 6015
rect 8128 5234 8156 6122
rect 8312 5710 8340 6598
rect 8300 5704 8352 5710
rect 8300 5646 8352 5652
rect 8404 5642 8432 6734
rect 8392 5636 8444 5642
rect 8392 5578 8444 5584
rect 8208 5568 8260 5574
rect 8208 5510 8260 5516
rect 8116 5228 8168 5234
rect 8116 5170 8168 5176
rect 8024 4616 8076 4622
rect 7748 4558 7800 4564
rect 7930 4584 7986 4593
rect 8024 4558 8076 4564
rect 8116 4616 8168 4622
rect 8116 4558 8168 4564
rect 7930 4519 7986 4528
rect 7610 4380 7918 4389
rect 7610 4378 7616 4380
rect 7672 4378 7696 4380
rect 7752 4378 7776 4380
rect 7832 4378 7856 4380
rect 7912 4378 7918 4380
rect 7672 4326 7674 4378
rect 7854 4326 7856 4378
rect 7610 4324 7616 4326
rect 7672 4324 7696 4326
rect 7752 4324 7776 4326
rect 7832 4324 7856 4326
rect 7912 4324 7918 4326
rect 7610 4315 7918 4324
rect 8128 4264 8156 4558
rect 8036 4236 8156 4264
rect 7472 4140 7524 4146
rect 7472 4082 7524 4088
rect 6920 3528 6972 3534
rect 6920 3470 6972 3476
rect 7012 3528 7064 3534
rect 7012 3470 7064 3476
rect 7380 3528 7432 3534
rect 7380 3470 7432 3476
rect 7484 3380 7512 4082
rect 8036 3398 8064 4236
rect 8220 4196 8248 5510
rect 8390 5400 8446 5409
rect 8390 5335 8446 5344
rect 8404 5098 8432 5335
rect 8392 5092 8444 5098
rect 8392 5034 8444 5040
rect 8300 5024 8352 5030
rect 8300 4966 8352 4972
rect 8312 4214 8340 4966
rect 8390 4448 8446 4457
rect 8390 4383 8446 4392
rect 8128 4168 8248 4196
rect 8300 4208 8352 4214
rect 8128 3602 8156 4168
rect 8300 4150 8352 4156
rect 8312 3942 8340 4150
rect 8404 4049 8432 4383
rect 8390 4040 8446 4049
rect 8390 3975 8446 3984
rect 8300 3936 8352 3942
rect 8300 3878 8352 3884
rect 8206 3632 8262 3641
rect 8116 3596 8168 3602
rect 8206 3567 8262 3576
rect 8116 3538 8168 3544
rect 8220 3534 8248 3567
rect 8208 3528 8260 3534
rect 8208 3470 8260 3476
rect 8300 3528 8352 3534
rect 8300 3470 8352 3476
rect 7286 3360 7342 3369
rect 7286 3295 7342 3304
rect 7392 3352 7512 3380
rect 8024 3392 8076 3398
rect 6736 3188 6788 3194
rect 6736 3130 6788 3136
rect 6552 3052 6604 3058
rect 6552 2994 6604 3000
rect 6644 3052 6696 3058
rect 6644 2994 6696 3000
rect 6460 2984 6512 2990
rect 6460 2926 6512 2932
rect 6472 1698 6500 2926
rect 6564 2854 6592 2994
rect 6644 2916 6696 2922
rect 6644 2858 6696 2864
rect 6736 2916 6788 2922
rect 6736 2858 6788 2864
rect 6552 2848 6604 2854
rect 6552 2790 6604 2796
rect 6550 2680 6606 2689
rect 6550 2615 6606 2624
rect 6564 2582 6592 2615
rect 6552 2576 6604 2582
rect 6552 2518 6604 2524
rect 6552 2440 6604 2446
rect 6552 2382 6604 2388
rect 6460 1692 6512 1698
rect 6460 1634 6512 1640
rect 6564 1601 6592 2382
rect 6550 1592 6606 1601
rect 6550 1527 6606 1536
rect 6368 1148 6420 1154
rect 6368 1090 6420 1096
rect 6000 876 6052 882
rect 6000 818 6052 824
rect 5264 672 5316 678
rect 5264 614 5316 620
rect 6656 610 6684 2858
rect 6748 2514 6776 2858
rect 6950 2748 7258 2757
rect 6950 2746 6956 2748
rect 7012 2746 7036 2748
rect 7092 2746 7116 2748
rect 7172 2746 7196 2748
rect 7252 2746 7258 2748
rect 7012 2694 7014 2746
rect 7194 2694 7196 2746
rect 6950 2692 6956 2694
rect 7012 2692 7036 2694
rect 7092 2692 7116 2694
rect 7172 2692 7196 2694
rect 7252 2692 7258 2694
rect 6950 2683 7258 2692
rect 6736 2508 6788 2514
rect 6736 2450 6788 2456
rect 6748 2106 6776 2450
rect 7196 2304 7248 2310
rect 7196 2246 7248 2252
rect 6736 2100 6788 2106
rect 6736 2042 6788 2048
rect 7208 1465 7236 2246
rect 7194 1456 7250 1465
rect 7194 1391 7250 1400
rect 7300 1222 7328 3295
rect 7288 1216 7340 1222
rect 7288 1158 7340 1164
rect 7392 1057 7420 3352
rect 8024 3334 8076 3340
rect 8208 3392 8260 3398
rect 8208 3334 8260 3340
rect 7610 3292 7918 3301
rect 7610 3290 7616 3292
rect 7672 3290 7696 3292
rect 7752 3290 7776 3292
rect 7832 3290 7856 3292
rect 7912 3290 7918 3292
rect 7672 3238 7674 3290
rect 7854 3238 7856 3290
rect 7610 3236 7616 3238
rect 7672 3236 7696 3238
rect 7752 3236 7776 3238
rect 7832 3236 7856 3238
rect 7912 3236 7918 3238
rect 7610 3227 7918 3236
rect 7472 3188 7524 3194
rect 7472 3130 7524 3136
rect 7484 2514 7512 3130
rect 7656 3120 7708 3126
rect 7656 3062 7708 3068
rect 7472 2508 7524 2514
rect 7472 2450 7524 2456
rect 7668 2310 7696 3062
rect 7932 2984 7984 2990
rect 7930 2952 7932 2961
rect 7984 2952 7986 2961
rect 8220 2922 8248 3334
rect 8312 3233 8340 3470
rect 8298 3224 8354 3233
rect 8298 3159 8354 3168
rect 8404 3080 8432 3975
rect 8496 3466 8524 10662
rect 8574 10568 8630 10577
rect 8574 10503 8630 10512
rect 8588 9042 8616 10503
rect 8576 9036 8628 9042
rect 8576 8978 8628 8984
rect 8680 8634 8708 12124
rect 8760 12106 8812 12112
rect 8760 11212 8812 11218
rect 8760 11154 8812 11160
rect 8668 8628 8720 8634
rect 8668 8570 8720 8576
rect 8576 8492 8628 8498
rect 8576 8434 8628 8440
rect 8668 8492 8720 8498
rect 8668 8434 8720 8440
rect 8588 8362 8616 8434
rect 8576 8356 8628 8362
rect 8576 8298 8628 8304
rect 8588 6458 8616 8298
rect 8680 7528 8708 8434
rect 8772 8294 8800 11154
rect 8760 8288 8812 8294
rect 8760 8230 8812 8236
rect 8864 7546 8892 14742
rect 8956 13938 8984 15399
rect 9128 14476 9180 14482
rect 9128 14418 9180 14424
rect 8944 13932 8996 13938
rect 8944 13874 8996 13880
rect 9140 13870 9168 14418
rect 9232 14074 9260 16050
rect 9508 15706 9536 17274
rect 9784 17270 9812 17478
rect 9772 17264 9824 17270
rect 9772 17206 9824 17212
rect 9588 17128 9640 17134
rect 9588 17070 9640 17076
rect 9312 15700 9364 15706
rect 9312 15642 9364 15648
rect 9496 15700 9548 15706
rect 9496 15642 9548 15648
rect 9324 15502 9352 15642
rect 9312 15496 9364 15502
rect 9312 15438 9364 15444
rect 9404 15428 9456 15434
rect 9404 15370 9456 15376
rect 9312 14952 9364 14958
rect 9312 14894 9364 14900
rect 9324 14482 9352 14894
rect 9312 14476 9364 14482
rect 9312 14418 9364 14424
rect 9310 14376 9366 14385
rect 9310 14311 9366 14320
rect 9324 14074 9352 14311
rect 9220 14068 9272 14074
rect 9220 14010 9272 14016
rect 9312 14068 9364 14074
rect 9312 14010 9364 14016
rect 9312 13932 9364 13938
rect 9312 13874 9364 13880
rect 9128 13864 9180 13870
rect 9128 13806 9180 13812
rect 9220 13864 9272 13870
rect 9220 13806 9272 13812
rect 9036 13524 9088 13530
rect 9036 13466 9088 13472
rect 9048 12782 9076 13466
rect 9036 12776 9088 12782
rect 9036 12718 9088 12724
rect 9036 12436 9088 12442
rect 9036 12378 9088 12384
rect 8944 12368 8996 12374
rect 8944 12310 8996 12316
rect 8956 11626 8984 12310
rect 8944 11620 8996 11626
rect 8944 11562 8996 11568
rect 8944 11076 8996 11082
rect 8944 11018 8996 11024
rect 8956 10062 8984 11018
rect 8944 10056 8996 10062
rect 8944 9998 8996 10004
rect 8944 9920 8996 9926
rect 8944 9862 8996 9868
rect 8852 7540 8904 7546
rect 8680 7500 8800 7528
rect 8668 7404 8720 7410
rect 8668 7346 8720 7352
rect 8680 6474 8708 7346
rect 8772 7002 8800 7500
rect 8852 7482 8904 7488
rect 8852 7336 8904 7342
rect 8852 7278 8904 7284
rect 8760 6996 8812 7002
rect 8760 6938 8812 6944
rect 8772 6662 8800 6938
rect 8864 6866 8892 7278
rect 8956 6934 8984 9862
rect 9048 9722 9076 12378
rect 9036 9716 9088 9722
rect 9036 9658 9088 9664
rect 9036 9580 9088 9586
rect 9036 9522 9088 9528
rect 9048 9353 9076 9522
rect 9034 9344 9090 9353
rect 9034 9279 9090 9288
rect 9036 9036 9088 9042
rect 9036 8978 9088 8984
rect 8944 6928 8996 6934
rect 8944 6870 8996 6876
rect 8852 6860 8904 6866
rect 8852 6802 8904 6808
rect 8956 6746 8984 6870
rect 9048 6769 9076 8978
rect 9140 7886 9168 13806
rect 9232 13297 9260 13806
rect 9324 13394 9352 13874
rect 9312 13388 9364 13394
rect 9312 13330 9364 13336
rect 9218 13288 9274 13297
rect 9218 13223 9274 13232
rect 9310 13152 9366 13161
rect 9310 13087 9366 13096
rect 9220 12980 9272 12986
rect 9220 12922 9272 12928
rect 9232 12238 9260 12922
rect 9324 12850 9352 13087
rect 9312 12844 9364 12850
rect 9312 12786 9364 12792
rect 9220 12232 9272 12238
rect 9220 12174 9272 12180
rect 9232 11393 9260 12174
rect 9312 12164 9364 12170
rect 9312 12106 9364 12112
rect 9218 11384 9274 11393
rect 9218 11319 9274 11328
rect 9220 11076 9272 11082
rect 9220 11018 9272 11024
rect 9232 9042 9260 11018
rect 9220 9036 9272 9042
rect 9220 8978 9272 8984
rect 9218 8936 9274 8945
rect 9218 8871 9274 8880
rect 9128 7880 9180 7886
rect 9128 7822 9180 7828
rect 8864 6718 8984 6746
rect 9034 6760 9090 6769
rect 8760 6656 8812 6662
rect 8760 6598 8812 6604
rect 8576 6452 8628 6458
rect 8680 6446 8800 6474
rect 8576 6394 8628 6400
rect 8588 4622 8616 6394
rect 8668 5092 8720 5098
rect 8668 5034 8720 5040
rect 8576 4616 8628 4622
rect 8576 4558 8628 4564
rect 8574 3904 8630 3913
rect 8574 3839 8630 3848
rect 8484 3460 8536 3466
rect 8484 3402 8536 3408
rect 8392 3074 8444 3080
rect 8300 3052 8352 3058
rect 8392 3016 8444 3022
rect 8300 2994 8352 3000
rect 8312 2961 8340 2994
rect 8588 2990 8616 3839
rect 8576 2984 8628 2990
rect 8298 2952 8354 2961
rect 7930 2887 7986 2896
rect 8208 2916 8260 2922
rect 8298 2887 8354 2896
rect 8404 2944 8576 2972
rect 8208 2858 8260 2864
rect 7840 2848 7892 2854
rect 7840 2790 7892 2796
rect 7852 2394 7880 2790
rect 8206 2680 8262 2689
rect 8206 2615 8262 2624
rect 7852 2366 7972 2394
rect 8220 2378 8248 2615
rect 7656 2304 7708 2310
rect 7470 2272 7526 2281
rect 7656 2246 7708 2252
rect 7944 2258 7972 2366
rect 8208 2372 8260 2378
rect 8208 2314 8260 2320
rect 8022 2272 8078 2281
rect 7944 2230 8022 2258
rect 7470 2207 7526 2216
rect 7484 1766 7512 2207
rect 7610 2204 7918 2213
rect 8022 2207 8078 2216
rect 7610 2202 7616 2204
rect 7672 2202 7696 2204
rect 7752 2202 7776 2204
rect 7832 2202 7856 2204
rect 7912 2202 7918 2204
rect 7672 2150 7674 2202
rect 7854 2150 7856 2202
rect 7610 2148 7616 2150
rect 7672 2148 7696 2150
rect 7752 2148 7776 2150
rect 7832 2148 7856 2150
rect 7912 2148 7918 2150
rect 7610 2139 7918 2148
rect 7472 1760 7524 1766
rect 7472 1702 7524 1708
rect 8404 1193 8432 2944
rect 8576 2926 8628 2932
rect 8680 2774 8708 5034
rect 8772 4672 8800 6446
rect 8864 5914 8892 6718
rect 9034 6695 9090 6704
rect 8942 6624 8998 6633
rect 8942 6559 8998 6568
rect 8956 6118 8984 6559
rect 8944 6112 8996 6118
rect 8944 6054 8996 6060
rect 8942 5944 8998 5953
rect 8852 5908 8904 5914
rect 8942 5879 8944 5888
rect 8852 5850 8904 5856
rect 8996 5879 8998 5888
rect 8944 5850 8996 5856
rect 8944 5704 8996 5710
rect 8944 5646 8996 5652
rect 8852 5296 8904 5302
rect 8850 5264 8852 5273
rect 8904 5264 8906 5273
rect 8850 5199 8906 5208
rect 8956 5166 8984 5646
rect 9048 5234 9076 6695
rect 9140 5846 9168 7822
rect 9128 5840 9180 5846
rect 9128 5782 9180 5788
rect 9128 5704 9180 5710
rect 9128 5646 9180 5652
rect 9140 5574 9168 5646
rect 9128 5568 9180 5574
rect 9126 5536 9128 5545
rect 9180 5536 9182 5545
rect 9126 5471 9182 5480
rect 9036 5228 9088 5234
rect 9036 5170 9088 5176
rect 9128 5228 9180 5234
rect 9128 5170 9180 5176
rect 8944 5160 8996 5166
rect 8944 5102 8996 5108
rect 9140 4758 9168 5170
rect 9128 4752 9180 4758
rect 9128 4694 9180 4700
rect 8772 4644 8984 4672
rect 8852 4548 8904 4554
rect 8852 4490 8904 4496
rect 8760 4480 8812 4486
rect 8864 4457 8892 4490
rect 8760 4422 8812 4428
rect 8850 4448 8906 4457
rect 8772 4214 8800 4422
rect 8850 4383 8906 4392
rect 8760 4208 8812 4214
rect 8760 4150 8812 4156
rect 8772 3466 8800 4150
rect 8850 4040 8906 4049
rect 8850 3975 8906 3984
rect 8760 3460 8812 3466
rect 8760 3402 8812 3408
rect 8496 2746 8708 2774
rect 8496 2514 8524 2746
rect 8666 2680 8722 2689
rect 8666 2615 8722 2624
rect 8574 2544 8630 2553
rect 8484 2508 8536 2514
rect 8680 2514 8708 2615
rect 8574 2479 8576 2488
rect 8484 2450 8536 2456
rect 8628 2479 8630 2488
rect 8668 2508 8720 2514
rect 8576 2450 8628 2456
rect 8668 2450 8720 2456
rect 8772 2446 8800 3402
rect 8864 3398 8892 3975
rect 8956 3913 8984 4644
rect 8942 3904 8998 3913
rect 8942 3839 8998 3848
rect 8852 3392 8904 3398
rect 8852 3334 8904 3340
rect 8956 3194 8984 3839
rect 9232 3534 9260 8871
rect 9324 8498 9352 12106
rect 9312 8492 9364 8498
rect 9312 8434 9364 8440
rect 9416 8294 9444 15370
rect 9496 14816 9548 14822
rect 9496 14758 9548 14764
rect 9508 14618 9536 14758
rect 9496 14612 9548 14618
rect 9496 14554 9548 14560
rect 9600 13870 9628 17070
rect 9862 16552 9918 16561
rect 9862 16487 9918 16496
rect 9772 15360 9824 15366
rect 9772 15302 9824 15308
rect 9784 15162 9812 15302
rect 9772 15156 9824 15162
rect 9772 15098 9824 15104
rect 9770 15056 9826 15065
rect 9770 14991 9772 15000
rect 9824 14991 9826 15000
rect 9772 14962 9824 14968
rect 9680 14952 9732 14958
rect 9680 14894 9732 14900
rect 9588 13864 9640 13870
rect 9588 13806 9640 13812
rect 9496 13524 9548 13530
rect 9496 13466 9548 13472
rect 9508 11880 9536 13466
rect 9692 12889 9720 14894
rect 9770 14376 9826 14385
rect 9770 14311 9826 14320
rect 9784 14278 9812 14311
rect 9772 14272 9824 14278
rect 9772 14214 9824 14220
rect 9876 13394 9904 16487
rect 10048 15972 10100 15978
rect 10048 15914 10100 15920
rect 9956 15156 10008 15162
rect 9956 15098 10008 15104
rect 9864 13388 9916 13394
rect 9864 13330 9916 13336
rect 9864 13252 9916 13258
rect 9864 13194 9916 13200
rect 9876 13025 9904 13194
rect 9862 13016 9918 13025
rect 9862 12951 9918 12960
rect 9678 12880 9734 12889
rect 9968 12832 9996 15098
rect 10060 13530 10088 15914
rect 10244 15026 10272 18566
rect 10874 18527 10930 18536
rect 10784 18012 10836 18018
rect 10784 17954 10836 17960
rect 10508 17128 10560 17134
rect 10508 17070 10560 17076
rect 10416 17060 10468 17066
rect 10416 17002 10468 17008
rect 10428 16590 10456 17002
rect 10520 16726 10548 17070
rect 10796 16726 10824 17954
rect 10508 16720 10560 16726
rect 10508 16662 10560 16668
rect 10692 16720 10744 16726
rect 10692 16662 10744 16668
rect 10784 16720 10836 16726
rect 10784 16662 10836 16668
rect 10416 16584 10468 16590
rect 10416 16526 10468 16532
rect 10600 16584 10652 16590
rect 10600 16526 10652 16532
rect 10508 16448 10560 16454
rect 10508 16390 10560 16396
rect 10416 16040 10468 16046
rect 10416 15982 10468 15988
rect 10324 15904 10376 15910
rect 10324 15846 10376 15852
rect 10140 15020 10192 15026
rect 10140 14962 10192 14968
rect 10232 15020 10284 15026
rect 10232 14962 10284 14968
rect 10048 13524 10100 13530
rect 10048 13466 10100 13472
rect 10060 12850 10088 13466
rect 10152 13433 10180 14962
rect 10232 13456 10284 13462
rect 10138 13424 10194 13433
rect 10232 13398 10284 13404
rect 10138 13359 10194 13368
rect 10138 12880 10194 12889
rect 9678 12815 9734 12824
rect 9876 12804 9996 12832
rect 10048 12844 10100 12850
rect 9772 12776 9824 12782
rect 9770 12744 9772 12753
rect 9824 12744 9826 12753
rect 9588 12708 9640 12714
rect 9770 12679 9826 12688
rect 9588 12650 9640 12656
rect 9600 12170 9628 12650
rect 9772 12436 9824 12442
rect 9876 12434 9904 12804
rect 10138 12815 10194 12824
rect 10048 12786 10100 12792
rect 9956 12708 10008 12714
rect 9956 12650 10008 12656
rect 9968 12617 9996 12650
rect 10152 12628 10180 12815
rect 9954 12608 10010 12617
rect 9954 12543 10010 12552
rect 10060 12600 10180 12628
rect 9824 12406 9904 12434
rect 9772 12378 9824 12384
rect 9680 12368 9732 12374
rect 10060 12356 10088 12600
rect 10140 12436 10192 12442
rect 10140 12378 10192 12384
rect 9680 12310 9732 12316
rect 9876 12328 10088 12356
rect 9588 12164 9640 12170
rect 9588 12106 9640 12112
rect 9692 12073 9720 12310
rect 9772 12096 9824 12102
rect 9678 12064 9734 12073
rect 9772 12038 9824 12044
rect 9678 11999 9734 12008
rect 9784 11898 9812 12038
rect 9772 11892 9824 11898
rect 9508 11852 9628 11880
rect 9496 11756 9548 11762
rect 9496 11698 9548 11704
rect 9508 11218 9536 11698
rect 9496 11212 9548 11218
rect 9496 11154 9548 11160
rect 9496 11008 9548 11014
rect 9496 10950 9548 10956
rect 9508 10742 9536 10950
rect 9496 10736 9548 10742
rect 9496 10678 9548 10684
rect 9494 10296 9550 10305
rect 9600 10282 9628 11852
rect 9772 11834 9824 11840
rect 9680 11756 9732 11762
rect 9680 11698 9732 11704
rect 9692 11529 9720 11698
rect 9770 11656 9826 11665
rect 9770 11591 9826 11600
rect 9678 11520 9734 11529
rect 9678 11455 9734 11464
rect 9678 11248 9734 11257
rect 9678 11183 9734 11192
rect 9550 10254 9628 10282
rect 9494 10231 9550 10240
rect 9508 10130 9536 10231
rect 9496 10124 9548 10130
rect 9496 10066 9548 10072
rect 9496 9988 9548 9994
rect 9496 9930 9548 9936
rect 9508 9897 9536 9930
rect 9494 9888 9550 9897
rect 9494 9823 9550 9832
rect 9496 9580 9548 9586
rect 9496 9522 9548 9528
rect 9312 8288 9364 8294
rect 9312 8230 9364 8236
rect 9404 8288 9456 8294
rect 9404 8230 9456 8236
rect 9324 7886 9352 8230
rect 9312 7880 9364 7886
rect 9312 7822 9364 7828
rect 9310 7168 9366 7177
rect 9310 7103 9366 7112
rect 9324 3534 9352 7103
rect 9416 4214 9444 8230
rect 9508 7800 9536 9522
rect 9588 9444 9640 9450
rect 9588 9386 9640 9392
rect 9600 8498 9628 9386
rect 9588 8492 9640 8498
rect 9588 8434 9640 8440
rect 9692 8378 9720 11183
rect 9784 10985 9812 11591
rect 9770 10976 9826 10985
rect 9770 10911 9826 10920
rect 9772 10736 9824 10742
rect 9772 10678 9824 10684
rect 9784 9518 9812 10678
rect 9772 9512 9824 9518
rect 9876 9489 9904 12328
rect 9954 12200 10010 12209
rect 9954 12135 10010 12144
rect 9968 11694 9996 12135
rect 10152 12050 10180 12378
rect 10244 12238 10272 13398
rect 10336 12374 10364 15846
rect 10428 15502 10456 15982
rect 10416 15496 10468 15502
rect 10416 15438 10468 15444
rect 10520 15065 10548 16390
rect 10612 16289 10640 16526
rect 10598 16280 10654 16289
rect 10598 16215 10654 16224
rect 10704 15978 10732 16662
rect 10888 16454 10916 18527
rect 11164 17202 11192 19200
rect 11520 18828 11572 18834
rect 11520 18770 11572 18776
rect 11532 18426 11560 18770
rect 11428 18420 11480 18426
rect 11428 18362 11480 18368
rect 11520 18420 11572 18426
rect 11520 18362 11572 18368
rect 11440 18222 11468 18362
rect 11428 18216 11480 18222
rect 11428 18158 11480 18164
rect 12346 17912 12402 17921
rect 12346 17847 12402 17856
rect 11152 17196 11204 17202
rect 11152 17138 11204 17144
rect 11980 17128 12032 17134
rect 11808 17088 11980 17116
rect 11336 16992 11388 16998
rect 11336 16934 11388 16940
rect 11518 16960 11574 16969
rect 11348 16697 11376 16934
rect 11518 16895 11574 16904
rect 11334 16688 11390 16697
rect 11334 16623 11390 16632
rect 11532 16522 11560 16895
rect 11612 16584 11664 16590
rect 11612 16526 11664 16532
rect 11336 16516 11388 16522
rect 11336 16458 11388 16464
rect 11520 16516 11572 16522
rect 11520 16458 11572 16464
rect 10876 16448 10928 16454
rect 10876 16390 10928 16396
rect 10888 16130 10916 16390
rect 10796 16102 10916 16130
rect 10692 15972 10744 15978
rect 10692 15914 10744 15920
rect 10598 15736 10654 15745
rect 10598 15671 10600 15680
rect 10652 15671 10654 15680
rect 10692 15700 10744 15706
rect 10600 15642 10652 15648
rect 10692 15642 10744 15648
rect 10600 15496 10652 15502
rect 10598 15464 10600 15473
rect 10652 15464 10654 15473
rect 10598 15399 10654 15408
rect 10506 15056 10562 15065
rect 10506 14991 10562 15000
rect 10416 14952 10468 14958
rect 10416 14894 10468 14900
rect 10428 13841 10456 14894
rect 10520 14346 10548 14991
rect 10600 14816 10652 14822
rect 10600 14758 10652 14764
rect 10508 14340 10560 14346
rect 10508 14282 10560 14288
rect 10506 13968 10562 13977
rect 10506 13903 10562 13912
rect 10414 13832 10470 13841
rect 10414 13767 10470 13776
rect 10416 13728 10468 13734
rect 10416 13670 10468 13676
rect 10428 12918 10456 13670
rect 10416 12912 10468 12918
rect 10416 12854 10468 12860
rect 10416 12776 10468 12782
rect 10416 12718 10468 12724
rect 10324 12368 10376 12374
rect 10324 12310 10376 12316
rect 10232 12232 10284 12238
rect 10232 12174 10284 12180
rect 10152 12022 10272 12050
rect 10140 11892 10192 11898
rect 10140 11834 10192 11840
rect 10048 11824 10100 11830
rect 10048 11766 10100 11772
rect 9956 11688 10008 11694
rect 9956 11630 10008 11636
rect 10060 11626 10088 11766
rect 10048 11620 10100 11626
rect 10048 11562 10100 11568
rect 9954 11520 10010 11529
rect 9954 11455 10010 11464
rect 9968 10849 9996 11455
rect 10048 11144 10100 11150
rect 10048 11086 10100 11092
rect 10060 11014 10088 11086
rect 10048 11008 10100 11014
rect 10048 10950 10100 10956
rect 9954 10840 10010 10849
rect 9954 10775 10010 10784
rect 9956 10736 10008 10742
rect 9956 10678 10008 10684
rect 9772 9454 9824 9460
rect 9862 9480 9918 9489
rect 9784 9178 9812 9454
rect 9862 9415 9918 9424
rect 9772 9172 9824 9178
rect 9772 9114 9824 9120
rect 9770 8800 9826 8809
rect 9770 8735 9826 8744
rect 9784 8537 9812 8735
rect 9770 8528 9826 8537
rect 9770 8463 9826 8472
rect 9600 8350 9720 8378
rect 9772 8424 9824 8430
rect 9772 8366 9824 8372
rect 9600 8129 9628 8350
rect 9680 8288 9732 8294
rect 9784 8265 9812 8366
rect 9680 8230 9732 8236
rect 9770 8256 9826 8265
rect 9586 8120 9642 8129
rect 9586 8055 9642 8064
rect 9692 7868 9720 8230
rect 9770 8191 9826 8200
rect 9772 7880 9824 7886
rect 9692 7840 9772 7868
rect 9772 7822 9824 7828
rect 9508 7772 9628 7800
rect 9494 7712 9550 7721
rect 9494 7647 9550 7656
rect 9508 6866 9536 7647
rect 9600 7546 9628 7772
rect 9678 7712 9734 7721
rect 9678 7647 9734 7656
rect 9588 7540 9640 7546
rect 9588 7482 9640 7488
rect 9692 7410 9720 7647
rect 9772 7540 9824 7546
rect 9772 7482 9824 7488
rect 9680 7404 9732 7410
rect 9680 7346 9732 7352
rect 9496 6860 9548 6866
rect 9496 6802 9548 6808
rect 9586 6760 9642 6769
rect 9586 6695 9642 6704
rect 9600 6497 9628 6695
rect 9680 6656 9732 6662
rect 9680 6598 9732 6604
rect 9586 6488 9642 6497
rect 9692 6458 9720 6598
rect 9586 6423 9642 6432
rect 9680 6452 9732 6458
rect 9496 6248 9548 6254
rect 9496 6190 9548 6196
rect 9508 5817 9536 6190
rect 9494 5808 9550 5817
rect 9494 5743 9550 5752
rect 9404 4208 9456 4214
rect 9600 4162 9628 6423
rect 9680 6394 9732 6400
rect 9678 6352 9734 6361
rect 9678 6287 9680 6296
rect 9732 6287 9734 6296
rect 9680 6258 9732 6264
rect 9784 5642 9812 7482
rect 9876 7410 9904 9415
rect 9968 8906 9996 10678
rect 10048 10056 10100 10062
rect 10048 9998 10100 10004
rect 9956 8900 10008 8906
rect 9956 8842 10008 8848
rect 10060 8786 10088 9998
rect 10152 8974 10180 11834
rect 10244 10305 10272 12022
rect 10336 11218 10364 12310
rect 10324 11212 10376 11218
rect 10324 11154 10376 11160
rect 10230 10296 10286 10305
rect 10230 10231 10286 10240
rect 10428 10180 10456 12718
rect 10520 12646 10548 13903
rect 10612 12889 10640 14758
rect 10704 14618 10732 15642
rect 10692 14612 10744 14618
rect 10692 14554 10744 14560
rect 10692 14408 10744 14414
rect 10692 14350 10744 14356
rect 10598 12880 10654 12889
rect 10598 12815 10654 12824
rect 10704 12730 10732 14350
rect 10796 13025 10824 16102
rect 10876 16040 10928 16046
rect 10876 15982 10928 15988
rect 10888 14793 10916 15982
rect 11152 15632 11204 15638
rect 11152 15574 11204 15580
rect 11060 15496 11112 15502
rect 11060 15438 11112 15444
rect 10968 15360 11020 15366
rect 10968 15302 11020 15308
rect 10874 14784 10930 14793
rect 10874 14719 10930 14728
rect 10888 13394 10916 14719
rect 10980 14618 11008 15302
rect 10968 14612 11020 14618
rect 10968 14554 11020 14560
rect 10966 14512 11022 14521
rect 10966 14447 11022 14456
rect 10980 14278 11008 14447
rect 10968 14272 11020 14278
rect 10968 14214 11020 14220
rect 10968 13864 11020 13870
rect 10968 13806 11020 13812
rect 10876 13388 10928 13394
rect 10876 13330 10928 13336
rect 10980 13138 11008 13806
rect 11072 13462 11100 15438
rect 11164 14890 11192 15574
rect 11244 15088 11296 15094
rect 11244 15030 11296 15036
rect 11152 14884 11204 14890
rect 11152 14826 11204 14832
rect 11256 14657 11284 15030
rect 11242 14648 11298 14657
rect 11242 14583 11298 14592
rect 11152 14544 11204 14550
rect 11152 14486 11204 14492
rect 11244 14544 11296 14550
rect 11244 14486 11296 14492
rect 11164 14074 11192 14486
rect 11152 14068 11204 14074
rect 11152 14010 11204 14016
rect 11060 13456 11112 13462
rect 11060 13398 11112 13404
rect 10980 13110 11100 13138
rect 10782 13016 10838 13025
rect 10782 12951 10838 12960
rect 11072 12889 11100 13110
rect 10874 12880 10930 12889
rect 11058 12880 11114 12889
rect 10874 12815 10876 12824
rect 10928 12815 10930 12824
rect 10968 12844 11020 12850
rect 10876 12786 10928 12792
rect 11058 12815 11114 12824
rect 10968 12786 11020 12792
rect 10600 12708 10652 12714
rect 10704 12702 10824 12730
rect 10600 12650 10652 12656
rect 10508 12640 10560 12646
rect 10508 12582 10560 12588
rect 10520 11880 10548 12582
rect 10612 12481 10640 12650
rect 10692 12640 10744 12646
rect 10692 12582 10744 12588
rect 10598 12472 10654 12481
rect 10598 12407 10654 12416
rect 10704 12238 10732 12582
rect 10692 12232 10744 12238
rect 10692 12174 10744 12180
rect 10520 11852 10640 11880
rect 10508 11756 10560 11762
rect 10508 11698 10560 11704
rect 10244 10152 10456 10180
rect 10140 8968 10192 8974
rect 10140 8910 10192 8916
rect 9968 8758 10088 8786
rect 9968 8294 9996 8758
rect 10046 8664 10102 8673
rect 10152 8634 10180 8910
rect 10046 8599 10102 8608
rect 10140 8628 10192 8634
rect 9956 8288 10008 8294
rect 9956 8230 10008 8236
rect 9954 8120 10010 8129
rect 9954 8055 10010 8064
rect 9968 7954 9996 8055
rect 9956 7948 10008 7954
rect 9956 7890 10008 7896
rect 9864 7404 9916 7410
rect 9864 7346 9916 7352
rect 9956 7336 10008 7342
rect 9956 7278 10008 7284
rect 9968 6914 9996 7278
rect 9876 6886 9996 6914
rect 9876 6633 9904 6886
rect 9862 6624 9918 6633
rect 9862 6559 9918 6568
rect 9772 5636 9824 5642
rect 9772 5578 9824 5584
rect 9680 4752 9732 4758
rect 9680 4694 9732 4700
rect 9692 4593 9720 4694
rect 9678 4584 9734 4593
rect 9678 4519 9734 4528
rect 9404 4150 9456 4156
rect 9508 4134 9628 4162
rect 9678 4176 9734 4185
rect 9404 3936 9456 3942
rect 9404 3878 9456 3884
rect 9220 3528 9272 3534
rect 9220 3470 9272 3476
rect 9312 3528 9364 3534
rect 9312 3470 9364 3476
rect 8944 3188 8996 3194
rect 8944 3130 8996 3136
rect 9128 3120 9180 3126
rect 9128 3062 9180 3068
rect 8852 2984 8904 2990
rect 8852 2926 8904 2932
rect 8864 2825 8892 2926
rect 8850 2816 8906 2825
rect 8850 2751 8906 2760
rect 9034 2680 9090 2689
rect 9034 2615 9036 2624
rect 9088 2615 9090 2624
rect 9036 2586 9088 2592
rect 8760 2440 8812 2446
rect 8482 2408 8538 2417
rect 8760 2382 8812 2388
rect 8482 2343 8538 2352
rect 8496 1562 8524 2343
rect 9140 2310 9168 3062
rect 9312 3052 9364 3058
rect 9312 2994 9364 3000
rect 9220 2644 9272 2650
rect 9220 2586 9272 2592
rect 9232 2446 9260 2586
rect 9324 2582 9352 2994
rect 9312 2576 9364 2582
rect 9312 2518 9364 2524
rect 9416 2514 9444 3878
rect 9508 3534 9536 4134
rect 9678 4111 9734 4120
rect 9588 4072 9640 4078
rect 9586 4040 9588 4049
rect 9640 4040 9642 4049
rect 9586 3975 9642 3984
rect 9692 3738 9720 4111
rect 9772 4072 9824 4078
rect 9772 4014 9824 4020
rect 9680 3732 9732 3738
rect 9680 3674 9732 3680
rect 9680 3596 9732 3602
rect 9680 3538 9732 3544
rect 9496 3528 9548 3534
rect 9496 3470 9548 3476
rect 9494 3224 9550 3233
rect 9692 3210 9720 3538
rect 9550 3182 9720 3210
rect 9494 3159 9550 3168
rect 9588 3052 9640 3058
rect 9588 2994 9640 3000
rect 9404 2508 9456 2514
rect 9404 2450 9456 2456
rect 9220 2440 9272 2446
rect 9220 2382 9272 2388
rect 9312 2440 9364 2446
rect 9312 2382 9364 2388
rect 9128 2304 9180 2310
rect 9128 2246 9180 2252
rect 9232 2038 9260 2382
rect 9220 2032 9272 2038
rect 9220 1974 9272 1980
rect 9324 1902 9352 2382
rect 9416 2106 9444 2450
rect 9600 2446 9628 2994
rect 9588 2440 9640 2446
rect 9588 2382 9640 2388
rect 9404 2100 9456 2106
rect 9404 2042 9456 2048
rect 9312 1896 9364 1902
rect 9312 1838 9364 1844
rect 9784 1630 9812 4014
rect 9876 3466 9904 6559
rect 9954 6488 10010 6497
rect 9954 6423 10010 6432
rect 9968 5710 9996 6423
rect 10060 6390 10088 8599
rect 10140 8570 10192 8576
rect 10244 8514 10272 10152
rect 10520 10112 10548 11698
rect 10428 10084 10548 10112
rect 10324 9580 10376 9586
rect 10324 9522 10376 9528
rect 10336 9042 10364 9522
rect 10324 9036 10376 9042
rect 10324 8978 10376 8984
rect 10324 8900 10376 8906
rect 10324 8842 10376 8848
rect 10152 8486 10272 8514
rect 10336 8498 10364 8842
rect 10428 8838 10456 10084
rect 10612 9586 10640 11852
rect 10600 9580 10652 9586
rect 10600 9522 10652 9528
rect 10704 9382 10732 12174
rect 10796 12102 10824 12702
rect 10784 12096 10836 12102
rect 10784 12038 10836 12044
rect 10796 11762 10824 12038
rect 10876 11824 10928 11830
rect 10874 11792 10876 11801
rect 10928 11792 10930 11801
rect 10784 11756 10836 11762
rect 10874 11727 10930 11736
rect 10784 11698 10836 11704
rect 10980 11642 11008 12786
rect 11164 12646 11192 14010
rect 11256 13326 11284 14486
rect 11348 13410 11376 16458
rect 11624 16046 11652 16526
rect 11808 16425 11836 17088
rect 11980 17070 12032 17076
rect 12360 16969 12388 17847
rect 12610 17436 12918 17445
rect 12610 17434 12616 17436
rect 12672 17434 12696 17436
rect 12752 17434 12776 17436
rect 12832 17434 12856 17436
rect 12912 17434 12918 17436
rect 12672 17382 12674 17434
rect 12854 17382 12856 17434
rect 12610 17380 12616 17382
rect 12672 17380 12696 17382
rect 12752 17380 12776 17382
rect 12832 17380 12856 17382
rect 12912 17380 12918 17382
rect 12438 17368 12494 17377
rect 12610 17371 12918 17380
rect 12438 17303 12494 17312
rect 12346 16960 12402 16969
rect 11950 16892 12258 16901
rect 12346 16895 12402 16904
rect 11950 16890 11956 16892
rect 12012 16890 12036 16892
rect 12092 16890 12116 16892
rect 12172 16890 12196 16892
rect 12252 16890 12258 16892
rect 12012 16838 12014 16890
rect 12194 16838 12196 16890
rect 11950 16836 11956 16838
rect 12012 16836 12036 16838
rect 12092 16836 12116 16838
rect 12172 16836 12196 16838
rect 12252 16836 12258 16838
rect 11950 16827 12258 16836
rect 12452 16833 12480 17303
rect 13176 17264 13228 17270
rect 13176 17206 13228 17212
rect 12992 16992 13044 16998
rect 12992 16934 13044 16940
rect 12438 16824 12494 16833
rect 12438 16759 12494 16768
rect 12440 16652 12492 16658
rect 12440 16594 12492 16600
rect 11794 16416 11850 16425
rect 11794 16351 11850 16360
rect 12452 16164 12480 16594
rect 12610 16348 12918 16357
rect 12610 16346 12616 16348
rect 12672 16346 12696 16348
rect 12752 16346 12776 16348
rect 12832 16346 12856 16348
rect 12912 16346 12918 16348
rect 12672 16294 12674 16346
rect 12854 16294 12856 16346
rect 12610 16292 12616 16294
rect 12672 16292 12696 16294
rect 12752 16292 12776 16294
rect 12832 16292 12856 16294
rect 12912 16292 12918 16294
rect 12610 16283 12918 16292
rect 13004 16250 13032 16934
rect 12992 16244 13044 16250
rect 12992 16186 13044 16192
rect 12532 16176 12584 16182
rect 12254 16144 12310 16153
rect 12452 16136 12532 16164
rect 12310 16102 12388 16130
rect 12254 16079 12310 16088
rect 11612 16040 11664 16046
rect 11612 15982 11664 15988
rect 11612 15904 11664 15910
rect 11612 15846 11664 15852
rect 11520 15564 11572 15570
rect 11520 15506 11572 15512
rect 11428 15496 11480 15502
rect 11428 15438 11480 15444
rect 11440 15201 11468 15438
rect 11532 15366 11560 15506
rect 11520 15360 11572 15366
rect 11520 15302 11572 15308
rect 11426 15192 11482 15201
rect 11426 15127 11482 15136
rect 11520 14816 11572 14822
rect 11520 14758 11572 14764
rect 11532 14521 11560 14758
rect 11518 14512 11574 14521
rect 11518 14447 11574 14456
rect 11520 14272 11572 14278
rect 11520 14214 11572 14220
rect 11426 13832 11482 13841
rect 11426 13767 11482 13776
rect 11440 13734 11468 13767
rect 11428 13728 11480 13734
rect 11428 13670 11480 13676
rect 11348 13382 11468 13410
rect 11244 13320 11296 13326
rect 11242 13288 11244 13297
rect 11296 13288 11298 13297
rect 11242 13223 11298 13232
rect 11242 13016 11298 13025
rect 11242 12951 11298 12960
rect 11256 12850 11284 12951
rect 11244 12844 11296 12850
rect 11244 12786 11296 12792
rect 11336 12844 11388 12850
rect 11336 12786 11388 12792
rect 11348 12753 11376 12786
rect 11334 12744 11390 12753
rect 11334 12679 11390 12688
rect 11152 12640 11204 12646
rect 11152 12582 11204 12588
rect 11244 12640 11296 12646
rect 11244 12582 11296 12588
rect 11256 12374 11284 12582
rect 11244 12368 11296 12374
rect 11244 12310 11296 12316
rect 11336 12368 11388 12374
rect 11336 12310 11388 12316
rect 11060 11824 11112 11830
rect 11060 11766 11112 11772
rect 10888 11614 11008 11642
rect 10888 11354 10916 11614
rect 10966 11384 11022 11393
rect 10876 11348 10928 11354
rect 11072 11370 11100 11766
rect 11152 11756 11204 11762
rect 11152 11698 11204 11704
rect 11022 11342 11100 11370
rect 10966 11319 11022 11328
rect 10876 11290 10928 11296
rect 10784 11280 10836 11286
rect 10784 11222 10836 11228
rect 10966 11248 11022 11257
rect 10796 10470 10824 11222
rect 10966 11183 11022 11192
rect 10980 11150 11008 11183
rect 10968 11144 11020 11150
rect 10968 11086 11020 11092
rect 10980 10849 11008 11086
rect 10966 10840 11022 10849
rect 10966 10775 11022 10784
rect 10966 10704 11022 10713
rect 10966 10639 11022 10648
rect 11060 10668 11112 10674
rect 10980 10470 11008 10639
rect 11060 10610 11112 10616
rect 10784 10464 10836 10470
rect 10968 10464 11020 10470
rect 10784 10406 10836 10412
rect 10888 10424 10968 10452
rect 10784 9580 10836 9586
rect 10784 9522 10836 9528
rect 10600 9376 10652 9382
rect 10600 9318 10652 9324
rect 10692 9376 10744 9382
rect 10692 9318 10744 9324
rect 10506 9072 10562 9081
rect 10506 9007 10562 9016
rect 10416 8832 10468 8838
rect 10416 8774 10468 8780
rect 10428 8537 10456 8774
rect 10414 8528 10470 8537
rect 10324 8492 10376 8498
rect 10048 6384 10100 6390
rect 10048 6326 10100 6332
rect 10152 5914 10180 8486
rect 10414 8463 10470 8472
rect 10324 8434 10376 8440
rect 10232 8424 10284 8430
rect 10232 8366 10284 8372
rect 10244 7410 10272 8366
rect 10232 7404 10284 7410
rect 10232 7346 10284 7352
rect 10232 6384 10284 6390
rect 10232 6326 10284 6332
rect 10140 5908 10192 5914
rect 10140 5850 10192 5856
rect 9956 5704 10008 5710
rect 9956 5646 10008 5652
rect 10048 5092 10100 5098
rect 10048 5034 10100 5040
rect 9956 4820 10008 4826
rect 9956 4762 10008 4768
rect 9968 4554 9996 4762
rect 9956 4548 10008 4554
rect 9956 4490 10008 4496
rect 9956 4208 10008 4214
rect 9956 4150 10008 4156
rect 9864 3460 9916 3466
rect 9864 3402 9916 3408
rect 9876 2961 9904 3402
rect 9968 3126 9996 4150
rect 10060 4078 10088 5034
rect 10048 4072 10100 4078
rect 10048 4014 10100 4020
rect 10244 3738 10272 6326
rect 10232 3732 10284 3738
rect 10232 3674 10284 3680
rect 9956 3120 10008 3126
rect 9956 3062 10008 3068
rect 9862 2952 9918 2961
rect 9862 2887 9918 2896
rect 9956 2372 10008 2378
rect 9956 2314 10008 2320
rect 9772 1624 9824 1630
rect 9772 1566 9824 1572
rect 8484 1556 8536 1562
rect 8484 1498 8536 1504
rect 8390 1184 8446 1193
rect 8390 1119 8446 1128
rect 7378 1048 7434 1057
rect 7378 983 7434 992
rect 9968 800 9996 2314
rect 10336 1737 10364 8434
rect 10416 8356 10468 8362
rect 10416 8298 10468 8304
rect 10428 5302 10456 8298
rect 10520 5914 10548 9007
rect 10612 8362 10640 9318
rect 10796 9217 10824 9522
rect 10888 9518 10916 10424
rect 10968 10406 11020 10412
rect 11072 9897 11100 10610
rect 11058 9888 11114 9897
rect 11058 9823 11114 9832
rect 10968 9716 11020 9722
rect 10968 9658 11020 9664
rect 11060 9716 11112 9722
rect 11060 9658 11112 9664
rect 10876 9512 10928 9518
rect 10876 9454 10928 9460
rect 10980 9450 11008 9658
rect 10968 9444 11020 9450
rect 10968 9386 11020 9392
rect 10782 9208 10838 9217
rect 10692 9172 10744 9178
rect 10782 9143 10838 9152
rect 10692 9114 10744 9120
rect 10704 8634 10732 9114
rect 10876 9104 10928 9110
rect 10876 9046 10928 9052
rect 10966 9072 11022 9081
rect 10692 8628 10744 8634
rect 10692 8570 10744 8576
rect 10782 8528 10838 8537
rect 10782 8463 10838 8472
rect 10600 8356 10652 8362
rect 10600 8298 10652 8304
rect 10692 8288 10744 8294
rect 10692 8230 10744 8236
rect 10704 7954 10732 8230
rect 10692 7948 10744 7954
rect 10692 7890 10744 7896
rect 10796 7886 10824 8463
rect 10784 7880 10836 7886
rect 10784 7822 10836 7828
rect 10784 7744 10836 7750
rect 10784 7686 10836 7692
rect 10600 7540 10652 7546
rect 10600 7482 10652 7488
rect 10612 7342 10640 7482
rect 10796 7410 10824 7686
rect 10888 7546 10916 9046
rect 10966 9007 11022 9016
rect 10980 8498 11008 9007
rect 10968 8492 11020 8498
rect 10968 8434 11020 8440
rect 10876 7540 10928 7546
rect 10876 7482 10928 7488
rect 10784 7404 10836 7410
rect 10784 7346 10836 7352
rect 10600 7336 10652 7342
rect 10600 7278 10652 7284
rect 10600 7200 10652 7206
rect 10600 7142 10652 7148
rect 10508 5908 10560 5914
rect 10508 5850 10560 5856
rect 10612 5710 10640 7142
rect 10782 7032 10838 7041
rect 10782 6967 10838 6976
rect 10796 6662 10824 6967
rect 10980 6882 11008 8434
rect 11072 7478 11100 9658
rect 11164 8294 11192 11698
rect 11348 11336 11376 12310
rect 11440 11626 11468 13382
rect 11532 12986 11560 14214
rect 11624 13870 11652 15846
rect 11950 15804 12258 15813
rect 11950 15802 11956 15804
rect 12012 15802 12036 15804
rect 12092 15802 12116 15804
rect 12172 15802 12196 15804
rect 12252 15802 12258 15804
rect 12012 15750 12014 15802
rect 12194 15750 12196 15802
rect 11950 15748 11956 15750
rect 12012 15748 12036 15750
rect 12092 15748 12116 15750
rect 12172 15748 12196 15750
rect 12252 15748 12258 15750
rect 11950 15739 12258 15748
rect 12360 15745 12388 16102
rect 12346 15736 12402 15745
rect 12346 15671 12402 15680
rect 11704 15496 11756 15502
rect 11756 15456 11836 15484
rect 11704 15438 11756 15444
rect 11702 15192 11758 15201
rect 11702 15127 11758 15136
rect 11716 14822 11744 15127
rect 11704 14816 11756 14822
rect 11704 14758 11756 14764
rect 11716 14550 11744 14758
rect 11704 14544 11756 14550
rect 11704 14486 11756 14492
rect 11612 13864 11664 13870
rect 11612 13806 11664 13812
rect 11704 13864 11756 13870
rect 11704 13806 11756 13812
rect 11624 13274 11652 13806
rect 11716 13569 11744 13806
rect 11702 13560 11758 13569
rect 11702 13495 11758 13504
rect 11624 13246 11744 13274
rect 11808 13258 11836 15456
rect 12348 15428 12400 15434
rect 12348 15370 12400 15376
rect 11950 14716 12258 14725
rect 11950 14714 11956 14716
rect 12012 14714 12036 14716
rect 12092 14714 12116 14716
rect 12172 14714 12196 14716
rect 12252 14714 12258 14716
rect 12012 14662 12014 14714
rect 12194 14662 12196 14714
rect 11950 14660 11956 14662
rect 12012 14660 12036 14662
rect 12092 14660 12116 14662
rect 12172 14660 12196 14662
rect 12252 14660 12258 14662
rect 11950 14651 12258 14660
rect 11888 14612 11940 14618
rect 12256 14612 12308 14618
rect 11940 14572 12020 14600
rect 11888 14554 11940 14560
rect 11888 14340 11940 14346
rect 11888 14282 11940 14288
rect 11900 13977 11928 14282
rect 11992 14278 12020 14572
rect 12256 14554 12308 14560
rect 12070 14512 12126 14521
rect 12070 14447 12126 14456
rect 11980 14272 12032 14278
rect 12084 14249 12112 14447
rect 11980 14214 12032 14220
rect 12070 14240 12126 14249
rect 12070 14175 12126 14184
rect 11886 13968 11942 13977
rect 11886 13903 11942 13912
rect 12268 13734 12296 14554
rect 12256 13728 12308 13734
rect 12256 13670 12308 13676
rect 11950 13628 12258 13637
rect 11950 13626 11956 13628
rect 12012 13626 12036 13628
rect 12092 13626 12116 13628
rect 12172 13626 12196 13628
rect 12252 13626 12258 13628
rect 12012 13574 12014 13626
rect 12194 13574 12196 13626
rect 11950 13572 11956 13574
rect 12012 13572 12036 13574
rect 12092 13572 12116 13574
rect 12172 13572 12196 13574
rect 12252 13572 12258 13574
rect 11950 13563 12258 13572
rect 12360 13512 12388 15370
rect 12452 15026 12480 16136
rect 12532 16118 12584 16124
rect 13188 16130 13216 17206
rect 13648 17202 13676 19200
rect 14280 18760 14332 18766
rect 14280 18702 14332 18708
rect 13820 18148 13872 18154
rect 13820 18090 13872 18096
rect 13636 17196 13688 17202
rect 13636 17138 13688 17144
rect 13544 16788 13596 16794
rect 13544 16730 13596 16736
rect 13728 16788 13780 16794
rect 13728 16730 13780 16736
rect 13452 16516 13504 16522
rect 13452 16458 13504 16464
rect 12624 16108 12676 16114
rect 13188 16102 13308 16130
rect 12624 16050 12676 16056
rect 12532 15972 12584 15978
rect 12532 15914 12584 15920
rect 12440 15020 12492 15026
rect 12440 14962 12492 14968
rect 12452 14278 12480 14962
rect 12440 14272 12492 14278
rect 12440 14214 12492 14220
rect 12438 14104 12494 14113
rect 12438 14039 12494 14048
rect 12544 14056 12572 15914
rect 12636 15570 12664 16050
rect 12624 15564 12676 15570
rect 12624 15506 12676 15512
rect 12716 15564 12768 15570
rect 12716 15506 12768 15512
rect 12624 15428 12676 15434
rect 12728 15416 12756 15506
rect 12808 15496 12860 15502
rect 12676 15388 12756 15416
rect 12806 15464 12808 15473
rect 12860 15464 12862 15473
rect 12806 15399 12862 15408
rect 12992 15428 13044 15434
rect 12624 15370 12676 15376
rect 12992 15370 13044 15376
rect 12610 15260 12918 15269
rect 12610 15258 12616 15260
rect 12672 15258 12696 15260
rect 12752 15258 12776 15260
rect 12832 15258 12856 15260
rect 12912 15258 12918 15260
rect 12672 15206 12674 15258
rect 12854 15206 12856 15258
rect 12610 15204 12616 15206
rect 12672 15204 12696 15206
rect 12752 15204 12776 15206
rect 12832 15204 12856 15206
rect 12912 15204 12918 15206
rect 12610 15195 12918 15204
rect 12808 15088 12860 15094
rect 12808 15030 12860 15036
rect 12624 14884 12676 14890
rect 12624 14826 12676 14832
rect 12636 14618 12664 14826
rect 12820 14657 12848 15030
rect 12900 15020 12952 15026
rect 12900 14962 12952 14968
rect 12806 14648 12862 14657
rect 12624 14612 12676 14618
rect 12624 14554 12676 14560
rect 12716 14612 12768 14618
rect 12806 14583 12862 14592
rect 12716 14554 12768 14560
rect 12728 14414 12756 14554
rect 12716 14408 12768 14414
rect 12716 14350 12768 14356
rect 12912 14260 12940 14962
rect 13004 14793 13032 15370
rect 13084 14952 13136 14958
rect 13084 14894 13136 14900
rect 12990 14784 13046 14793
rect 12990 14719 13046 14728
rect 12992 14544 13044 14550
rect 12992 14486 13044 14492
rect 13004 14414 13032 14486
rect 12992 14408 13044 14414
rect 12992 14350 13044 14356
rect 12912 14232 13032 14260
rect 12610 14172 12918 14181
rect 12610 14170 12616 14172
rect 12672 14170 12696 14172
rect 12752 14170 12776 14172
rect 12832 14170 12856 14172
rect 12912 14170 12918 14172
rect 12672 14118 12674 14170
rect 12854 14118 12856 14170
rect 12610 14116 12616 14118
rect 12672 14116 12696 14118
rect 12752 14116 12776 14118
rect 12832 14116 12856 14118
rect 12912 14116 12918 14118
rect 12610 14107 12918 14116
rect 12452 13938 12480 14039
rect 12544 14028 12664 14056
rect 12440 13932 12492 13938
rect 12440 13874 12492 13880
rect 12440 13728 12492 13734
rect 12440 13670 12492 13676
rect 12532 13728 12584 13734
rect 12532 13670 12584 13676
rect 12084 13484 12388 13512
rect 11888 13388 11940 13394
rect 11888 13330 11940 13336
rect 11980 13388 12032 13394
rect 11980 13330 12032 13336
rect 11716 13190 11744 13246
rect 11796 13252 11848 13258
rect 11796 13194 11848 13200
rect 11612 13184 11664 13190
rect 11612 13126 11664 13132
rect 11704 13184 11756 13190
rect 11704 13126 11756 13132
rect 11520 12980 11572 12986
rect 11520 12922 11572 12928
rect 11624 12753 11652 13126
rect 11900 12986 11928 13330
rect 11888 12980 11940 12986
rect 11888 12922 11940 12928
rect 11702 12880 11758 12889
rect 11992 12850 12020 13330
rect 12084 12850 12112 13484
rect 12452 13394 12480 13670
rect 12440 13388 12492 13394
rect 12440 13330 12492 13336
rect 11702 12815 11758 12824
rect 11980 12844 12032 12850
rect 11716 12782 11744 12815
rect 11980 12786 12032 12792
rect 12072 12844 12124 12850
rect 12072 12786 12124 12792
rect 12440 12844 12492 12850
rect 12440 12786 12492 12792
rect 11704 12776 11756 12782
rect 11610 12744 11666 12753
rect 11704 12718 11756 12724
rect 11796 12776 11848 12782
rect 11796 12718 11848 12724
rect 12256 12776 12308 12782
rect 12308 12736 12388 12764
rect 12256 12718 12308 12724
rect 11610 12679 11666 12688
rect 11808 12628 11836 12718
rect 11518 12608 11574 12617
rect 11518 12543 11574 12552
rect 11716 12600 11836 12628
rect 11532 12434 11560 12543
rect 11532 12406 11652 12434
rect 11624 12306 11652 12406
rect 11612 12300 11664 12306
rect 11612 12242 11664 12248
rect 11520 11756 11572 11762
rect 11520 11698 11572 11704
rect 11428 11620 11480 11626
rect 11428 11562 11480 11568
rect 11348 11308 11468 11336
rect 11244 11212 11296 11218
rect 11244 11154 11296 11160
rect 11256 10577 11284 11154
rect 11440 11098 11468 11308
rect 11348 11070 11468 11098
rect 11242 10568 11298 10577
rect 11242 10503 11298 10512
rect 11256 9518 11284 10503
rect 11244 9512 11296 9518
rect 11244 9454 11296 9460
rect 11348 9178 11376 11070
rect 11532 10792 11560 11698
rect 11624 11014 11652 12242
rect 11716 11150 11744 12600
rect 11950 12540 12258 12549
rect 11950 12538 11956 12540
rect 12012 12538 12036 12540
rect 12092 12538 12116 12540
rect 12172 12538 12196 12540
rect 12252 12538 12258 12540
rect 12012 12486 12014 12538
rect 12194 12486 12196 12538
rect 11950 12484 11956 12486
rect 12012 12484 12036 12486
rect 12092 12484 12116 12486
rect 12172 12484 12196 12486
rect 12252 12484 12258 12486
rect 11794 12472 11850 12481
rect 11950 12475 12258 12484
rect 11794 12407 11850 12416
rect 11808 11801 11836 12407
rect 12256 12096 12308 12102
rect 12256 12038 12308 12044
rect 11794 11792 11850 11801
rect 11794 11727 11850 11736
rect 11796 11620 11848 11626
rect 11796 11562 11848 11568
rect 11704 11144 11756 11150
rect 11704 11086 11756 11092
rect 11612 11008 11664 11014
rect 11808 10962 11836 11562
rect 12268 11540 12296 12038
rect 12360 11694 12388 12736
rect 12452 12306 12480 12786
rect 12440 12300 12492 12306
rect 12440 12242 12492 12248
rect 12438 11928 12494 11937
rect 12438 11863 12494 11872
rect 12348 11688 12400 11694
rect 12348 11630 12400 11636
rect 12268 11512 12388 11540
rect 11950 11452 12258 11461
rect 11950 11450 11956 11452
rect 12012 11450 12036 11452
rect 12092 11450 12116 11452
rect 12172 11450 12196 11452
rect 12252 11450 12258 11452
rect 12012 11398 12014 11450
rect 12194 11398 12196 11450
rect 11950 11396 11956 11398
rect 12012 11396 12036 11398
rect 12092 11396 12116 11398
rect 12172 11396 12196 11398
rect 12252 11396 12258 11398
rect 11950 11387 12258 11396
rect 11888 11144 11940 11150
rect 11888 11086 11940 11092
rect 12070 11112 12126 11121
rect 11612 10950 11664 10956
rect 11440 10764 11560 10792
rect 11336 9172 11388 9178
rect 11336 9114 11388 9120
rect 11348 8566 11376 9114
rect 11336 8560 11388 8566
rect 11336 8502 11388 8508
rect 11336 8356 11388 8362
rect 11336 8298 11388 8304
rect 11152 8288 11204 8294
rect 11152 8230 11204 8236
rect 11244 8016 11296 8022
rect 11348 7993 11376 8298
rect 11244 7958 11296 7964
rect 11334 7984 11390 7993
rect 11152 7744 11204 7750
rect 11152 7686 11204 7692
rect 11060 7472 11112 7478
rect 11060 7414 11112 7420
rect 11072 7041 11100 7414
rect 11164 7206 11192 7686
rect 11152 7200 11204 7206
rect 11152 7142 11204 7148
rect 11058 7032 11114 7041
rect 11058 6967 11114 6976
rect 10980 6854 11192 6882
rect 10876 6792 10928 6798
rect 10876 6734 10928 6740
rect 11060 6792 11112 6798
rect 11060 6734 11112 6740
rect 10784 6656 10836 6662
rect 10784 6598 10836 6604
rect 10692 6316 10744 6322
rect 10692 6258 10744 6264
rect 10784 6316 10836 6322
rect 10784 6258 10836 6264
rect 10600 5704 10652 5710
rect 10520 5664 10600 5692
rect 10520 5302 10548 5664
rect 10600 5646 10652 5652
rect 10600 5568 10652 5574
rect 10600 5510 10652 5516
rect 10612 5370 10640 5510
rect 10600 5364 10652 5370
rect 10600 5306 10652 5312
rect 10416 5296 10468 5302
rect 10416 5238 10468 5244
rect 10508 5296 10560 5302
rect 10508 5238 10560 5244
rect 10428 4622 10456 5238
rect 10600 5024 10652 5030
rect 10600 4966 10652 4972
rect 10416 4616 10468 4622
rect 10416 4558 10468 4564
rect 10416 4072 10468 4078
rect 10416 4014 10468 4020
rect 10428 3194 10456 4014
rect 10416 3188 10468 3194
rect 10416 3130 10468 3136
rect 10612 2854 10640 4966
rect 10704 4622 10732 6258
rect 10796 5794 10824 6258
rect 10888 5914 10916 6734
rect 10968 6384 11020 6390
rect 10968 6326 11020 6332
rect 10876 5908 10928 5914
rect 10876 5850 10928 5856
rect 10796 5766 10916 5794
rect 10784 5568 10836 5574
rect 10888 5545 10916 5766
rect 10784 5510 10836 5516
rect 10874 5536 10930 5545
rect 10796 5001 10824 5510
rect 10874 5471 10930 5480
rect 10876 5364 10928 5370
rect 10876 5306 10928 5312
rect 10782 4992 10838 5001
rect 10782 4927 10838 4936
rect 10692 4616 10744 4622
rect 10692 4558 10744 4564
rect 10692 4480 10744 4486
rect 10692 4422 10744 4428
rect 10600 2848 10652 2854
rect 10600 2790 10652 2796
rect 10704 1970 10732 4422
rect 10888 3670 10916 5306
rect 10980 5234 11008 6326
rect 10968 5228 11020 5234
rect 10968 5170 11020 5176
rect 10968 4140 11020 4146
rect 10968 4082 11020 4088
rect 10980 4049 11008 4082
rect 10966 4040 11022 4049
rect 10966 3975 11022 3984
rect 10876 3664 10928 3670
rect 10876 3606 10928 3612
rect 10876 3460 10928 3466
rect 10876 3402 10928 3408
rect 10784 3052 10836 3058
rect 10784 2994 10836 3000
rect 10796 2961 10824 2994
rect 10782 2952 10838 2961
rect 10782 2887 10838 2896
rect 10784 2848 10836 2854
rect 10784 2790 10836 2796
rect 10796 2106 10824 2790
rect 10888 2446 10916 3402
rect 11072 3126 11100 6734
rect 11164 5710 11192 6854
rect 11256 6118 11284 7958
rect 11334 7919 11390 7928
rect 11336 7200 11388 7206
rect 11336 7142 11388 7148
rect 11244 6112 11296 6118
rect 11244 6054 11296 6060
rect 11152 5704 11204 5710
rect 11152 5646 11204 5652
rect 11164 4146 11192 5646
rect 11152 4140 11204 4146
rect 11152 4082 11204 4088
rect 11164 3942 11192 4082
rect 11152 3936 11204 3942
rect 11152 3878 11204 3884
rect 11256 3482 11284 6054
rect 11348 4078 11376 7142
rect 11336 4072 11388 4078
rect 11336 4014 11388 4020
rect 11440 4026 11468 10764
rect 11518 10704 11574 10713
rect 11624 10674 11652 10950
rect 11716 10934 11836 10962
rect 11518 10639 11520 10648
rect 11572 10639 11574 10648
rect 11612 10668 11664 10674
rect 11520 10610 11572 10616
rect 11612 10610 11664 10616
rect 11532 10538 11560 10610
rect 11520 10532 11572 10538
rect 11520 10474 11572 10480
rect 11520 10260 11572 10266
rect 11520 10202 11572 10208
rect 11532 7750 11560 10202
rect 11624 9178 11652 10610
rect 11716 9466 11744 10934
rect 11796 10804 11848 10810
rect 11796 10746 11848 10752
rect 11808 10674 11836 10746
rect 11900 10742 11928 11086
rect 11980 11076 12032 11082
rect 12070 11047 12126 11056
rect 11980 11018 12032 11024
rect 11888 10736 11940 10742
rect 11888 10678 11940 10684
rect 11796 10668 11848 10674
rect 11796 10610 11848 10616
rect 11808 10538 11836 10610
rect 11796 10532 11848 10538
rect 11796 10474 11848 10480
rect 11992 10452 12020 11018
rect 12084 10606 12112 11047
rect 12164 11008 12216 11014
rect 12360 10996 12388 11512
rect 12452 11393 12480 11863
rect 12438 11384 12494 11393
rect 12438 11319 12494 11328
rect 12544 11218 12572 13670
rect 12636 13326 12664 14028
rect 12716 13932 12768 13938
rect 12716 13874 12768 13880
rect 12728 13734 12756 13874
rect 12716 13728 12768 13734
rect 12716 13670 12768 13676
rect 12624 13320 12676 13326
rect 12624 13262 12676 13268
rect 12610 13084 12918 13093
rect 12610 13082 12616 13084
rect 12672 13082 12696 13084
rect 12752 13082 12776 13084
rect 12832 13082 12856 13084
rect 12912 13082 12918 13084
rect 12672 13030 12674 13082
rect 12854 13030 12856 13082
rect 12610 13028 12616 13030
rect 12672 13028 12696 13030
rect 12752 13028 12776 13030
rect 12832 13028 12856 13030
rect 12912 13028 12918 13030
rect 12610 13019 12918 13028
rect 12900 12844 12952 12850
rect 12900 12786 12952 12792
rect 12716 12776 12768 12782
rect 12716 12718 12768 12724
rect 12624 12640 12676 12646
rect 12624 12582 12676 12588
rect 12636 12238 12664 12582
rect 12624 12232 12676 12238
rect 12624 12174 12676 12180
rect 12728 12102 12756 12718
rect 12716 12096 12768 12102
rect 12912 12084 12940 12786
rect 13004 12442 13032 14232
rect 13096 13326 13124 14894
rect 13176 14884 13228 14890
rect 13176 14826 13228 14832
rect 13188 14113 13216 14826
rect 13174 14104 13230 14113
rect 13174 14039 13230 14048
rect 13176 13932 13228 13938
rect 13176 13874 13228 13880
rect 13084 13320 13136 13326
rect 13084 13262 13136 13268
rect 13082 13016 13138 13025
rect 13082 12951 13138 12960
rect 13096 12918 13124 12951
rect 13084 12912 13136 12918
rect 13084 12854 13136 12860
rect 13188 12714 13216 13874
rect 13280 13326 13308 16102
rect 13464 15026 13492 16458
rect 13556 16182 13584 16730
rect 13544 16176 13596 16182
rect 13544 16118 13596 16124
rect 13740 15094 13768 16730
rect 13728 15088 13780 15094
rect 13728 15030 13780 15036
rect 13832 15026 13860 18090
rect 13910 16960 13966 16969
rect 13910 16895 13966 16904
rect 13360 15020 13412 15026
rect 13360 14962 13412 14968
rect 13452 15020 13504 15026
rect 13452 14962 13504 14968
rect 13820 15020 13872 15026
rect 13820 14962 13872 14968
rect 13372 14929 13400 14962
rect 13358 14920 13414 14929
rect 13358 14855 13414 14864
rect 13360 14544 13412 14550
rect 13360 14486 13412 14492
rect 13636 14544 13688 14550
rect 13636 14486 13688 14492
rect 13268 13320 13320 13326
rect 13268 13262 13320 13268
rect 13268 12912 13320 12918
rect 13268 12854 13320 12860
rect 13176 12708 13228 12714
rect 13176 12650 13228 12656
rect 12992 12436 13044 12442
rect 12992 12378 13044 12384
rect 13084 12300 13136 12306
rect 13084 12242 13136 12248
rect 12992 12232 13044 12238
rect 12990 12200 12992 12209
rect 13044 12200 13046 12209
rect 12990 12135 13046 12144
rect 12912 12056 13032 12084
rect 12716 12038 12768 12044
rect 12610 11996 12918 12005
rect 12610 11994 12616 11996
rect 12672 11994 12696 11996
rect 12752 11994 12776 11996
rect 12832 11994 12856 11996
rect 12912 11994 12918 11996
rect 12672 11942 12674 11994
rect 12854 11942 12856 11994
rect 12610 11940 12616 11942
rect 12672 11940 12696 11942
rect 12752 11940 12776 11942
rect 12832 11940 12856 11942
rect 12912 11940 12918 11942
rect 12610 11931 12918 11940
rect 12808 11892 12860 11898
rect 12808 11834 12860 11840
rect 12820 11762 12848 11834
rect 12808 11756 12860 11762
rect 12808 11698 12860 11704
rect 12716 11280 12768 11286
rect 12716 11222 12768 11228
rect 12532 11212 12584 11218
rect 12532 11154 12584 11160
rect 12728 11150 12756 11222
rect 12716 11144 12768 11150
rect 12716 11086 12768 11092
rect 12440 11076 12492 11082
rect 12440 11018 12492 11024
rect 12216 10968 12388 10996
rect 12164 10950 12216 10956
rect 12176 10674 12204 10950
rect 12452 10849 12480 11018
rect 12610 10908 12918 10917
rect 12610 10906 12616 10908
rect 12672 10906 12696 10908
rect 12752 10906 12776 10908
rect 12832 10906 12856 10908
rect 12912 10906 12918 10908
rect 12672 10854 12674 10906
rect 12854 10854 12856 10906
rect 12610 10852 12616 10854
rect 12672 10852 12696 10854
rect 12752 10852 12776 10854
rect 12832 10852 12856 10854
rect 12912 10852 12918 10854
rect 12438 10840 12494 10849
rect 12610 10843 12918 10852
rect 12438 10775 12494 10784
rect 12624 10804 12676 10810
rect 12624 10746 12676 10752
rect 12164 10668 12216 10674
rect 12164 10610 12216 10616
rect 12072 10600 12124 10606
rect 12072 10542 12124 10548
rect 11992 10424 12388 10452
rect 11950 10364 12258 10373
rect 11950 10362 11956 10364
rect 12012 10362 12036 10364
rect 12092 10362 12116 10364
rect 12172 10362 12196 10364
rect 12252 10362 12258 10364
rect 12012 10310 12014 10362
rect 12194 10310 12196 10362
rect 11950 10308 11956 10310
rect 12012 10308 12036 10310
rect 12092 10308 12116 10310
rect 12172 10308 12196 10310
rect 12252 10308 12258 10310
rect 11794 10296 11850 10305
rect 11950 10299 12258 10308
rect 11850 10240 11928 10248
rect 11794 10231 11928 10240
rect 11808 10220 11928 10231
rect 11716 9438 11836 9466
rect 11704 9376 11756 9382
rect 11704 9318 11756 9324
rect 11612 9172 11664 9178
rect 11612 9114 11664 9120
rect 11610 9072 11666 9081
rect 11610 9007 11612 9016
rect 11664 9007 11666 9016
rect 11612 8978 11664 8984
rect 11520 7744 11572 7750
rect 11520 7686 11572 7692
rect 11610 7712 11666 7721
rect 11610 7647 11666 7656
rect 11520 7540 11572 7546
rect 11520 7482 11572 7488
rect 11532 7410 11560 7482
rect 11624 7410 11652 7647
rect 11520 7404 11572 7410
rect 11520 7346 11572 7352
rect 11612 7404 11664 7410
rect 11612 7346 11664 7352
rect 11532 5370 11560 7346
rect 11610 7168 11666 7177
rect 11610 7103 11666 7112
rect 11624 6798 11652 7103
rect 11612 6792 11664 6798
rect 11612 6734 11664 6740
rect 11716 6610 11744 9318
rect 11808 9160 11836 9438
rect 11900 9382 11928 10220
rect 12360 10112 12388 10424
rect 12532 10260 12584 10266
rect 12532 10202 12584 10208
rect 12176 10084 12388 10112
rect 12176 9874 12204 10084
rect 12254 10024 12310 10033
rect 12310 9982 12480 10010
rect 12254 9959 12310 9968
rect 12348 9920 12400 9926
rect 12176 9846 12296 9874
rect 12348 9862 12400 9868
rect 12162 9752 12218 9761
rect 12268 9722 12296 9846
rect 12162 9687 12164 9696
rect 12216 9687 12218 9696
rect 12256 9716 12308 9722
rect 12164 9658 12216 9664
rect 12256 9658 12308 9664
rect 12360 9654 12388 9862
rect 12348 9648 12400 9654
rect 12348 9590 12400 9596
rect 11888 9376 11940 9382
rect 11888 9318 11940 9324
rect 12348 9376 12400 9382
rect 12348 9318 12400 9324
rect 11950 9276 12258 9285
rect 11950 9274 11956 9276
rect 12012 9274 12036 9276
rect 12092 9274 12116 9276
rect 12172 9274 12196 9276
rect 12252 9274 12258 9276
rect 12012 9222 12014 9274
rect 12194 9222 12196 9274
rect 11950 9220 11956 9222
rect 12012 9220 12036 9222
rect 12092 9220 12116 9222
rect 12172 9220 12196 9222
rect 12252 9220 12258 9222
rect 11950 9211 12258 9220
rect 12164 9172 12216 9178
rect 11808 9132 12112 9160
rect 11888 8832 11940 8838
rect 11888 8774 11940 8780
rect 11900 8537 11928 8774
rect 11886 8528 11942 8537
rect 11886 8463 11942 8472
rect 12084 8276 12112 9132
rect 12164 9114 12216 9120
rect 12176 8566 12204 9114
rect 12254 8800 12310 8809
rect 12254 8735 12310 8744
rect 12164 8560 12216 8566
rect 12164 8502 12216 8508
rect 12268 8498 12296 8735
rect 12256 8492 12308 8498
rect 12256 8434 12308 8440
rect 11624 6582 11744 6610
rect 11808 8248 12112 8276
rect 11624 5692 11652 6582
rect 11704 6452 11756 6458
rect 11704 6394 11756 6400
rect 11716 6236 11744 6394
rect 11808 6390 11836 8248
rect 11950 8188 12258 8197
rect 11950 8186 11956 8188
rect 12012 8186 12036 8188
rect 12092 8186 12116 8188
rect 12172 8186 12196 8188
rect 12252 8186 12258 8188
rect 12012 8134 12014 8186
rect 12194 8134 12196 8186
rect 11950 8132 11956 8134
rect 12012 8132 12036 8134
rect 12092 8132 12116 8134
rect 12172 8132 12196 8134
rect 12252 8132 12258 8134
rect 11950 8123 12258 8132
rect 12360 8072 12388 9318
rect 12452 9178 12480 9982
rect 12544 9674 12572 10202
rect 12636 9926 12664 10746
rect 12716 10668 12768 10674
rect 12716 10610 12768 10616
rect 12900 10668 12952 10674
rect 12900 10610 12952 10616
rect 12728 10441 12756 10610
rect 12808 10600 12860 10606
rect 12808 10542 12860 10548
rect 12714 10432 12770 10441
rect 12714 10367 12770 10376
rect 12820 9926 12848 10542
rect 12624 9920 12676 9926
rect 12624 9862 12676 9868
rect 12808 9920 12860 9926
rect 12912 9908 12940 10610
rect 13004 10266 13032 12056
rect 13096 11132 13124 12242
rect 13176 12232 13228 12238
rect 13174 12200 13176 12209
rect 13228 12200 13230 12209
rect 13174 12135 13230 12144
rect 13176 12096 13228 12102
rect 13176 12038 13228 12044
rect 13188 11150 13216 12038
rect 13280 11626 13308 12854
rect 13372 12102 13400 14486
rect 13452 14476 13504 14482
rect 13452 14418 13504 14424
rect 13464 13841 13492 14418
rect 13544 14340 13596 14346
rect 13544 14282 13596 14288
rect 13450 13832 13506 13841
rect 13450 13767 13506 13776
rect 13452 13728 13504 13734
rect 13452 13670 13504 13676
rect 13464 12850 13492 13670
rect 13452 12844 13504 12850
rect 13452 12786 13504 12792
rect 13452 12708 13504 12714
rect 13452 12650 13504 12656
rect 13360 12096 13412 12102
rect 13360 12038 13412 12044
rect 13360 11892 13412 11898
rect 13360 11834 13412 11840
rect 13268 11620 13320 11626
rect 13268 11562 13320 11568
rect 13266 11520 13322 11529
rect 13266 11455 13322 11464
rect 13176 11144 13228 11150
rect 13096 11104 13146 11132
rect 13118 10724 13146 11104
rect 13176 11086 13228 11092
rect 13280 10996 13308 11455
rect 13096 10696 13146 10724
rect 13188 10968 13308 10996
rect 12992 10260 13044 10266
rect 12992 10202 13044 10208
rect 12912 9880 13032 9908
rect 12808 9862 12860 9868
rect 12610 9820 12918 9829
rect 12610 9818 12616 9820
rect 12672 9818 12696 9820
rect 12752 9818 12776 9820
rect 12832 9818 12856 9820
rect 12912 9818 12918 9820
rect 12672 9766 12674 9818
rect 12854 9766 12856 9818
rect 12610 9764 12616 9766
rect 12672 9764 12696 9766
rect 12752 9764 12776 9766
rect 12832 9764 12856 9766
rect 12912 9764 12918 9766
rect 12610 9755 12918 9764
rect 13004 9704 13032 9880
rect 12912 9676 13032 9704
rect 12544 9646 12664 9674
rect 12532 9580 12584 9586
rect 12532 9522 12584 9528
rect 12544 9450 12572 9522
rect 12532 9444 12584 9450
rect 12532 9386 12584 9392
rect 12440 9172 12492 9178
rect 12440 9114 12492 9120
rect 12530 9072 12586 9081
rect 12452 9030 12530 9058
rect 12452 8090 12480 9030
rect 12636 9042 12664 9646
rect 12808 9648 12860 9654
rect 12808 9590 12860 9596
rect 12530 9007 12586 9016
rect 12624 9036 12676 9042
rect 12624 8978 12676 8984
rect 12820 8974 12848 9590
rect 12808 8968 12860 8974
rect 12808 8910 12860 8916
rect 12532 8900 12584 8906
rect 12532 8842 12584 8848
rect 12268 8044 12388 8072
rect 12440 8084 12492 8090
rect 11978 7440 12034 7449
rect 11978 7375 11980 7384
rect 12032 7375 12034 7384
rect 11980 7346 12032 7352
rect 12268 7206 12296 8044
rect 12440 8026 12492 8032
rect 12348 7336 12400 7342
rect 12348 7278 12400 7284
rect 12256 7200 12308 7206
rect 12256 7142 12308 7148
rect 11950 7100 12258 7109
rect 11950 7098 11956 7100
rect 12012 7098 12036 7100
rect 12092 7098 12116 7100
rect 12172 7098 12196 7100
rect 12252 7098 12258 7100
rect 12012 7046 12014 7098
rect 12194 7046 12196 7098
rect 11950 7044 11956 7046
rect 12012 7044 12036 7046
rect 12092 7044 12116 7046
rect 12172 7044 12196 7046
rect 12252 7044 12258 7046
rect 11950 7035 12258 7044
rect 12256 6724 12308 6730
rect 12256 6666 12308 6672
rect 11796 6384 11848 6390
rect 11796 6326 11848 6332
rect 12268 6322 12296 6666
rect 12256 6316 12308 6322
rect 12256 6258 12308 6264
rect 11716 6208 11836 6236
rect 11808 5710 11836 6208
rect 11950 6012 12258 6021
rect 11950 6010 11956 6012
rect 12012 6010 12036 6012
rect 12092 6010 12116 6012
rect 12172 6010 12196 6012
rect 12252 6010 12258 6012
rect 12012 5958 12014 6010
rect 12194 5958 12196 6010
rect 11950 5956 11956 5958
rect 12012 5956 12036 5958
rect 12092 5956 12116 5958
rect 12172 5956 12196 5958
rect 12252 5956 12258 5958
rect 11950 5947 12258 5956
rect 11704 5704 11756 5710
rect 11624 5664 11704 5692
rect 11704 5646 11756 5652
rect 11796 5704 11848 5710
rect 11796 5646 11848 5652
rect 11612 5568 11664 5574
rect 11612 5510 11664 5516
rect 11520 5364 11572 5370
rect 11520 5306 11572 5312
rect 11518 5264 11574 5273
rect 11518 5199 11574 5208
rect 11532 4622 11560 5199
rect 11520 4616 11572 4622
rect 11520 4558 11572 4564
rect 11624 4468 11652 5510
rect 11716 4706 11744 5646
rect 11794 5536 11850 5545
rect 11794 5471 11850 5480
rect 11808 5166 11836 5471
rect 12254 5400 12310 5409
rect 12254 5335 12310 5344
rect 12268 5234 12296 5335
rect 12256 5228 12308 5234
rect 12256 5170 12308 5176
rect 11796 5160 11848 5166
rect 11796 5102 11848 5108
rect 12268 5030 12296 5170
rect 12256 5024 12308 5030
rect 12256 4966 12308 4972
rect 11950 4924 12258 4933
rect 11950 4922 11956 4924
rect 12012 4922 12036 4924
rect 12092 4922 12116 4924
rect 12172 4922 12196 4924
rect 12252 4922 12258 4924
rect 12012 4870 12014 4922
rect 12194 4870 12196 4922
rect 11950 4868 11956 4870
rect 12012 4868 12036 4870
rect 12092 4868 12116 4870
rect 12172 4868 12196 4870
rect 12252 4868 12258 4870
rect 11950 4859 12258 4868
rect 12072 4820 12124 4826
rect 12360 4808 12388 7278
rect 12544 6798 12572 8842
rect 12912 8838 12940 9676
rect 12992 9444 13044 9450
rect 12992 9386 13044 9392
rect 12900 8832 12952 8838
rect 12900 8774 12952 8780
rect 12610 8732 12918 8741
rect 12610 8730 12616 8732
rect 12672 8730 12696 8732
rect 12752 8730 12776 8732
rect 12832 8730 12856 8732
rect 12912 8730 12918 8732
rect 12672 8678 12674 8730
rect 12854 8678 12856 8730
rect 12610 8676 12616 8678
rect 12672 8676 12696 8678
rect 12752 8676 12776 8678
rect 12832 8676 12856 8678
rect 12912 8676 12918 8678
rect 12610 8667 12918 8676
rect 12808 8288 12860 8294
rect 13004 8265 13032 9386
rect 12808 8230 12860 8236
rect 12990 8256 13046 8265
rect 12622 8120 12678 8129
rect 12622 8055 12678 8064
rect 12636 7750 12664 8055
rect 12820 7750 12848 8230
rect 12990 8191 13046 8200
rect 12992 7948 13044 7954
rect 12992 7890 13044 7896
rect 12624 7744 12676 7750
rect 12624 7686 12676 7692
rect 12808 7744 12860 7750
rect 12808 7686 12860 7692
rect 12610 7644 12918 7653
rect 12610 7642 12616 7644
rect 12672 7642 12696 7644
rect 12752 7642 12776 7644
rect 12832 7642 12856 7644
rect 12912 7642 12918 7644
rect 12672 7590 12674 7642
rect 12854 7590 12856 7642
rect 12610 7588 12616 7590
rect 12672 7588 12696 7590
rect 12752 7588 12776 7590
rect 12832 7588 12856 7590
rect 12912 7588 12918 7590
rect 12610 7579 12918 7588
rect 13004 7274 13032 7890
rect 13096 7546 13124 10696
rect 13188 9602 13216 10968
rect 13266 10840 13322 10849
rect 13266 10775 13268 10784
rect 13320 10775 13322 10784
rect 13268 10746 13320 10752
rect 13268 10464 13320 10470
rect 13268 10406 13320 10412
rect 13280 10266 13308 10406
rect 13268 10260 13320 10266
rect 13268 10202 13320 10208
rect 13268 9988 13320 9994
rect 13268 9930 13320 9936
rect 13280 9761 13308 9930
rect 13266 9752 13322 9761
rect 13266 9687 13268 9696
rect 13320 9687 13322 9696
rect 13268 9658 13320 9664
rect 13188 9574 13308 9602
rect 13176 8628 13228 8634
rect 13176 8570 13228 8576
rect 13084 7540 13136 7546
rect 13084 7482 13136 7488
rect 12992 7268 13044 7274
rect 12992 7210 13044 7216
rect 12622 6896 12678 6905
rect 12622 6831 12678 6840
rect 12808 6860 12860 6866
rect 12636 6798 12664 6831
rect 12808 6802 12860 6808
rect 12992 6860 13044 6866
rect 12992 6802 13044 6808
rect 12532 6792 12584 6798
rect 12532 6734 12584 6740
rect 12624 6792 12676 6798
rect 12624 6734 12676 6740
rect 12820 6662 12848 6802
rect 12532 6656 12584 6662
rect 12532 6598 12584 6604
rect 12808 6656 12860 6662
rect 12808 6598 12860 6604
rect 12440 6248 12492 6254
rect 12440 6190 12492 6196
rect 12452 5953 12480 6190
rect 12544 6168 12572 6598
rect 12610 6556 12918 6565
rect 12610 6554 12616 6556
rect 12672 6554 12696 6556
rect 12752 6554 12776 6556
rect 12832 6554 12856 6556
rect 12912 6554 12918 6556
rect 12672 6502 12674 6554
rect 12854 6502 12856 6554
rect 12610 6500 12616 6502
rect 12672 6500 12696 6502
rect 12752 6500 12776 6502
rect 12832 6500 12856 6502
rect 12912 6500 12918 6502
rect 12610 6491 12918 6500
rect 12544 6140 12664 6168
rect 12438 5944 12494 5953
rect 12636 5914 12664 6140
rect 12714 6080 12770 6089
rect 12714 6015 12770 6024
rect 12438 5879 12494 5888
rect 12624 5908 12676 5914
rect 12624 5850 12676 5856
rect 12728 5534 12756 6015
rect 12544 5506 12756 5534
rect 12544 5302 12572 5506
rect 12610 5468 12918 5477
rect 12610 5466 12616 5468
rect 12672 5466 12696 5468
rect 12752 5466 12776 5468
rect 12832 5466 12856 5468
rect 12912 5466 12918 5468
rect 12672 5414 12674 5466
rect 12854 5414 12856 5466
rect 12610 5412 12616 5414
rect 12672 5412 12696 5414
rect 12752 5412 12776 5414
rect 12832 5412 12856 5414
rect 12912 5412 12918 5414
rect 12610 5403 12918 5412
rect 12532 5296 12584 5302
rect 12532 5238 12584 5244
rect 12532 5024 12584 5030
rect 12532 4966 12584 4972
rect 12124 4780 12388 4808
rect 12438 4856 12494 4865
rect 12438 4791 12494 4800
rect 12072 4762 12124 4768
rect 11716 4678 12020 4706
rect 11796 4616 11848 4622
rect 11794 4584 11796 4593
rect 11888 4616 11940 4622
rect 11848 4584 11850 4593
rect 11888 4558 11940 4564
rect 11794 4519 11850 4528
rect 11900 4468 11928 4558
rect 11624 4440 11928 4468
rect 11992 4214 12020 4678
rect 12452 4457 12480 4791
rect 12438 4448 12494 4457
rect 12438 4383 12494 4392
rect 12544 4264 12572 4966
rect 13004 4593 13032 6802
rect 13188 5710 13216 8570
rect 13176 5704 13228 5710
rect 13176 5646 13228 5652
rect 13084 5160 13136 5166
rect 13084 5102 13136 5108
rect 12990 4584 13046 4593
rect 12990 4519 13046 4528
rect 12610 4380 12918 4389
rect 12610 4378 12616 4380
rect 12672 4378 12696 4380
rect 12752 4378 12776 4380
rect 12832 4378 12856 4380
rect 12912 4378 12918 4380
rect 12672 4326 12674 4378
rect 12854 4326 12856 4378
rect 12610 4324 12616 4326
rect 12672 4324 12696 4326
rect 12752 4324 12776 4326
rect 12832 4324 12856 4326
rect 12912 4324 12918 4326
rect 12610 4315 12918 4324
rect 12992 4276 13044 4282
rect 12544 4236 12756 4264
rect 11980 4208 12032 4214
rect 11980 4150 12032 4156
rect 12346 4176 12402 4185
rect 12346 4111 12348 4120
rect 12400 4111 12402 4120
rect 12348 4082 12400 4088
rect 11796 4072 11848 4078
rect 11440 3998 11652 4026
rect 11796 4014 11848 4020
rect 11520 3936 11572 3942
rect 11520 3878 11572 3884
rect 11428 3732 11480 3738
rect 11428 3674 11480 3680
rect 11256 3454 11376 3482
rect 11060 3120 11112 3126
rect 11060 3062 11112 3068
rect 10968 3052 11020 3058
rect 10968 2994 11020 3000
rect 10876 2440 10928 2446
rect 10876 2382 10928 2388
rect 10784 2100 10836 2106
rect 10784 2042 10836 2048
rect 10980 2038 11008 2994
rect 11072 2514 11100 3062
rect 11244 2984 11296 2990
rect 11244 2926 11296 2932
rect 11060 2508 11112 2514
rect 11060 2450 11112 2456
rect 11152 2440 11204 2446
rect 11152 2382 11204 2388
rect 11060 2304 11112 2310
rect 11060 2246 11112 2252
rect 10968 2032 11020 2038
rect 10968 1974 11020 1980
rect 10692 1964 10744 1970
rect 10692 1906 10744 1912
rect 11072 1766 11100 2246
rect 11060 1760 11112 1766
rect 10322 1728 10378 1737
rect 11060 1702 11112 1708
rect 10322 1663 10378 1672
rect 11164 1358 11192 2382
rect 11152 1352 11204 1358
rect 11152 1294 11204 1300
rect 11256 1290 11284 2926
rect 11348 2854 11376 3454
rect 11336 2848 11388 2854
rect 11336 2790 11388 2796
rect 11440 2582 11468 3674
rect 11428 2576 11480 2582
rect 11428 2518 11480 2524
rect 11336 2440 11388 2446
rect 11334 2408 11336 2417
rect 11388 2408 11390 2417
rect 11334 2343 11390 2352
rect 11532 1834 11560 3878
rect 11624 3058 11652 3998
rect 11702 3904 11758 3913
rect 11702 3839 11758 3848
rect 11716 3738 11744 3839
rect 11704 3732 11756 3738
rect 11704 3674 11756 3680
rect 11702 3632 11758 3641
rect 11808 3602 11836 4014
rect 11950 3836 12258 3845
rect 11950 3834 11956 3836
rect 12012 3834 12036 3836
rect 12092 3834 12116 3836
rect 12172 3834 12196 3836
rect 12252 3834 12258 3836
rect 12012 3782 12014 3834
rect 12194 3782 12196 3834
rect 11950 3780 11956 3782
rect 12012 3780 12036 3782
rect 12092 3780 12116 3782
rect 12172 3780 12196 3782
rect 12252 3780 12258 3782
rect 11950 3771 12258 3780
rect 12346 3768 12402 3777
rect 12346 3703 12402 3712
rect 11702 3567 11758 3576
rect 11796 3596 11848 3602
rect 11716 3194 11744 3567
rect 11796 3538 11848 3544
rect 11704 3188 11756 3194
rect 11704 3130 11756 3136
rect 11612 3052 11664 3058
rect 11664 3012 11744 3040
rect 11612 2994 11664 3000
rect 11612 2848 11664 2854
rect 11612 2790 11664 2796
rect 11624 2446 11652 2790
rect 11716 2446 11744 3012
rect 11612 2440 11664 2446
rect 11612 2382 11664 2388
rect 11704 2440 11756 2446
rect 11704 2382 11756 2388
rect 11612 2304 11664 2310
rect 11612 2246 11664 2252
rect 11520 1828 11572 1834
rect 11520 1770 11572 1776
rect 11244 1284 11296 1290
rect 11244 1226 11296 1232
rect 6644 604 6696 610
rect 6644 546 6696 552
rect 3976 536 4028 542
rect 3882 504 3938 513
rect 3976 478 4028 484
rect 3882 439 3938 448
rect 9954 0 10010 800
rect 11624 649 11652 2246
rect 11808 1018 11836 3538
rect 11888 3528 11940 3534
rect 11888 3470 11940 3476
rect 11900 3126 11928 3470
rect 12072 3392 12124 3398
rect 12360 3369 12388 3703
rect 12728 3534 12756 4236
rect 12992 4218 13044 4224
rect 12808 3664 12860 3670
rect 12806 3632 12808 3641
rect 12860 3632 12862 3641
rect 12806 3567 12862 3576
rect 12624 3528 12676 3534
rect 12624 3470 12676 3476
rect 12716 3528 12768 3534
rect 12716 3470 12768 3476
rect 12636 3398 12664 3470
rect 12532 3392 12584 3398
rect 12072 3334 12124 3340
rect 12346 3360 12402 3369
rect 11888 3120 11940 3126
rect 11888 3062 11940 3068
rect 12084 3058 12112 3334
rect 12532 3334 12584 3340
rect 12624 3392 12676 3398
rect 12624 3334 12676 3340
rect 12346 3295 12402 3304
rect 12438 3224 12494 3233
rect 12438 3159 12494 3168
rect 12452 3058 12480 3159
rect 12072 3052 12124 3058
rect 12072 2994 12124 3000
rect 12440 3052 12492 3058
rect 12440 2994 12492 3000
rect 12348 2916 12400 2922
rect 12348 2858 12400 2864
rect 11950 2748 12258 2757
rect 11950 2746 11956 2748
rect 12012 2746 12036 2748
rect 12092 2746 12116 2748
rect 12172 2746 12196 2748
rect 12252 2746 12258 2748
rect 12012 2694 12014 2746
rect 12194 2694 12196 2746
rect 11950 2692 11956 2694
rect 12012 2692 12036 2694
rect 12092 2692 12116 2694
rect 12172 2692 12196 2694
rect 12252 2692 12258 2694
rect 11950 2683 12258 2692
rect 11978 2544 12034 2553
rect 11978 2479 12034 2488
rect 11992 2446 12020 2479
rect 11980 2440 12032 2446
rect 11980 2382 12032 2388
rect 11796 1012 11848 1018
rect 11796 954 11848 960
rect 12360 785 12388 2858
rect 12440 2440 12492 2446
rect 12440 2382 12492 2388
rect 12452 2310 12480 2382
rect 12440 2304 12492 2310
rect 12440 2246 12492 2252
rect 12346 776 12402 785
rect 12346 711 12402 720
rect 12544 678 12572 3334
rect 12610 3292 12918 3301
rect 12610 3290 12616 3292
rect 12672 3290 12696 3292
rect 12752 3290 12776 3292
rect 12832 3290 12856 3292
rect 12912 3290 12918 3292
rect 12672 3238 12674 3290
rect 12854 3238 12856 3290
rect 12610 3236 12616 3238
rect 12672 3236 12696 3238
rect 12752 3236 12776 3238
rect 12832 3236 12856 3238
rect 12912 3236 12918 3238
rect 12610 3227 12918 3236
rect 12716 2984 12768 2990
rect 13004 2972 13032 4218
rect 13096 4214 13124 5102
rect 13280 4554 13308 9574
rect 13372 8022 13400 11834
rect 13360 8016 13412 8022
rect 13360 7958 13412 7964
rect 13360 7744 13412 7750
rect 13360 7686 13412 7692
rect 13372 6322 13400 7686
rect 13464 7177 13492 12650
rect 13556 12646 13584 14282
rect 13648 14074 13676 14486
rect 13832 14226 13860 14962
rect 13924 14414 13952 16895
rect 14188 16516 14240 16522
rect 14188 16458 14240 16464
rect 14096 14612 14148 14618
rect 14096 14554 14148 14560
rect 13912 14408 13964 14414
rect 13912 14350 13964 14356
rect 13832 14198 13952 14226
rect 13636 14068 13688 14074
rect 13636 14010 13688 14016
rect 13820 14068 13872 14074
rect 13820 14010 13872 14016
rect 13728 13864 13780 13870
rect 13728 13806 13780 13812
rect 13636 13320 13688 13326
rect 13636 13262 13688 13268
rect 13544 12640 13596 12646
rect 13544 12582 13596 12588
rect 13556 12442 13584 12582
rect 13544 12436 13596 12442
rect 13544 12378 13596 12384
rect 13544 12300 13596 12306
rect 13544 12242 13596 12248
rect 13556 10690 13584 12242
rect 13648 10810 13676 13262
rect 13740 11830 13768 13806
rect 13728 11824 13780 11830
rect 13728 11766 13780 11772
rect 13728 11552 13780 11558
rect 13728 11494 13780 11500
rect 13636 10804 13688 10810
rect 13636 10746 13688 10752
rect 13556 10662 13676 10690
rect 13544 10600 13596 10606
rect 13544 10542 13596 10548
rect 13450 7168 13506 7177
rect 13450 7103 13506 7112
rect 13556 6934 13584 10542
rect 13648 9178 13676 10662
rect 13636 9172 13688 9178
rect 13636 9114 13688 9120
rect 13740 9110 13768 11494
rect 13832 11286 13860 14010
rect 13924 14006 13952 14198
rect 13912 14000 13964 14006
rect 13912 13942 13964 13948
rect 14004 13388 14056 13394
rect 14004 13330 14056 13336
rect 13912 12776 13964 12782
rect 13912 12718 13964 12724
rect 13924 11898 13952 12718
rect 14016 12170 14044 13330
rect 14004 12164 14056 12170
rect 14004 12106 14056 12112
rect 14002 11928 14058 11937
rect 13912 11892 13964 11898
rect 14002 11863 14058 11872
rect 13912 11834 13964 11840
rect 14016 11778 14044 11863
rect 13924 11750 14044 11778
rect 13924 11529 13952 11750
rect 14004 11688 14056 11694
rect 14004 11630 14056 11636
rect 13910 11520 13966 11529
rect 13910 11455 13966 11464
rect 13910 11384 13966 11393
rect 13910 11319 13966 11328
rect 13820 11280 13872 11286
rect 13820 11222 13872 11228
rect 13818 11112 13874 11121
rect 13818 11047 13874 11056
rect 13728 9104 13780 9110
rect 13728 9046 13780 9052
rect 13636 8968 13688 8974
rect 13636 8910 13688 8916
rect 13544 6928 13596 6934
rect 13544 6870 13596 6876
rect 13648 6712 13676 8910
rect 13728 8560 13780 8566
rect 13728 8502 13780 8508
rect 13740 8362 13768 8502
rect 13728 8356 13780 8362
rect 13728 8298 13780 8304
rect 13726 8256 13782 8265
rect 13726 8191 13782 8200
rect 13740 7818 13768 8191
rect 13832 7886 13860 11047
rect 13924 10470 13952 11319
rect 14016 10674 14044 11630
rect 14004 10668 14056 10674
rect 14004 10610 14056 10616
rect 14016 10538 14044 10610
rect 14004 10532 14056 10538
rect 14004 10474 14056 10480
rect 13912 10464 13964 10470
rect 13912 10406 13964 10412
rect 13924 9874 13952 10406
rect 13924 9846 14044 9874
rect 13912 9104 13964 9110
rect 13912 9046 13964 9052
rect 13924 8090 13952 9046
rect 14016 8974 14044 9846
rect 14004 8968 14056 8974
rect 14004 8910 14056 8916
rect 14004 8560 14056 8566
rect 14004 8502 14056 8508
rect 13912 8084 13964 8090
rect 13912 8026 13964 8032
rect 13910 7984 13966 7993
rect 13910 7919 13966 7928
rect 13924 7886 13952 7919
rect 13820 7880 13872 7886
rect 13820 7822 13872 7828
rect 13912 7880 13964 7886
rect 13912 7822 13964 7828
rect 13728 7812 13780 7818
rect 13728 7754 13780 7760
rect 13728 7268 13780 7274
rect 13728 7210 13780 7216
rect 13464 6684 13676 6712
rect 13360 6316 13412 6322
rect 13360 6258 13412 6264
rect 13268 4548 13320 4554
rect 13268 4490 13320 4496
rect 13084 4208 13136 4214
rect 13084 4150 13136 4156
rect 13372 3890 13400 6258
rect 13464 5234 13492 6684
rect 13634 6624 13690 6633
rect 13634 6559 13690 6568
rect 13544 5772 13596 5778
rect 13544 5714 13596 5720
rect 13452 5228 13504 5234
rect 13452 5170 13504 5176
rect 13464 4010 13492 5170
rect 13556 4622 13584 5714
rect 13648 4865 13676 6559
rect 13634 4856 13690 4865
rect 13634 4791 13690 4800
rect 13544 4616 13596 4622
rect 13596 4576 13676 4604
rect 13544 4558 13596 4564
rect 13542 4448 13598 4457
rect 13542 4383 13598 4392
rect 13452 4004 13504 4010
rect 13452 3946 13504 3952
rect 13280 3862 13400 3890
rect 13176 3664 13228 3670
rect 13176 3606 13228 3612
rect 13084 3052 13136 3058
rect 13084 2994 13136 3000
rect 12768 2944 13032 2972
rect 12716 2926 12768 2932
rect 12808 2440 12860 2446
rect 12860 2400 13032 2428
rect 12808 2382 12860 2388
rect 12610 2204 12918 2213
rect 12610 2202 12616 2204
rect 12672 2202 12696 2204
rect 12752 2202 12776 2204
rect 12832 2202 12856 2204
rect 12912 2202 12918 2204
rect 12672 2150 12674 2202
rect 12854 2150 12856 2202
rect 12610 2148 12616 2150
rect 12672 2148 12696 2150
rect 12752 2148 12776 2150
rect 12832 2148 12856 2150
rect 12912 2148 12918 2150
rect 12610 2139 12918 2148
rect 13004 1290 13032 2400
rect 13096 1494 13124 2994
rect 13188 2106 13216 3606
rect 13280 2310 13308 3862
rect 13464 3534 13492 3946
rect 13452 3528 13504 3534
rect 13452 3470 13504 3476
rect 13360 3392 13412 3398
rect 13360 3334 13412 3340
rect 13372 2922 13400 3334
rect 13360 2916 13412 2922
rect 13360 2858 13412 2864
rect 13372 2650 13400 2858
rect 13360 2644 13412 2650
rect 13360 2586 13412 2592
rect 13268 2304 13320 2310
rect 13268 2246 13320 2252
rect 13176 2100 13228 2106
rect 13176 2042 13228 2048
rect 13556 2038 13584 4383
rect 13648 3534 13676 4576
rect 13740 4078 13768 7210
rect 13728 4072 13780 4078
rect 13728 4014 13780 4020
rect 13636 3528 13688 3534
rect 13636 3470 13688 3476
rect 13648 3058 13676 3470
rect 13636 3052 13688 3058
rect 13636 2994 13688 3000
rect 13726 2680 13782 2689
rect 13726 2615 13782 2624
rect 13740 2446 13768 2615
rect 13832 2514 13860 7822
rect 13912 7268 13964 7274
rect 13912 7210 13964 7216
rect 13924 4146 13952 7210
rect 14016 6662 14044 8502
rect 14004 6656 14056 6662
rect 14004 6598 14056 6604
rect 14108 6458 14136 14554
rect 14200 14346 14228 16458
rect 14292 15094 14320 18702
rect 15936 18556 15988 18562
rect 15936 18498 15988 18504
rect 14464 18488 14516 18494
rect 14464 18430 14516 18436
rect 14372 18284 14424 18290
rect 14372 18226 14424 18232
rect 14280 15088 14332 15094
rect 14280 15030 14332 15036
rect 14278 14512 14334 14521
rect 14278 14447 14334 14456
rect 14292 14414 14320 14447
rect 14280 14408 14332 14414
rect 14280 14350 14332 14356
rect 14188 14340 14240 14346
rect 14188 14282 14240 14288
rect 14200 13433 14228 14282
rect 14384 14226 14412 18226
rect 14292 14198 14412 14226
rect 14186 13424 14242 13433
rect 14186 13359 14242 13368
rect 14188 12640 14240 12646
rect 14188 12582 14240 12588
rect 14200 12209 14228 12582
rect 14292 12345 14320 14198
rect 14476 14090 14504 18430
rect 14648 18352 14700 18358
rect 14648 18294 14700 18300
rect 14554 16688 14610 16697
rect 14554 16623 14610 16632
rect 14384 14062 14504 14090
rect 14278 12336 14334 12345
rect 14278 12271 14334 12280
rect 14186 12200 14242 12209
rect 14186 12135 14242 12144
rect 14280 12164 14332 12170
rect 14280 12106 14332 12112
rect 14292 12073 14320 12106
rect 14278 12064 14334 12073
rect 14278 11999 14334 12008
rect 14186 11384 14242 11393
rect 14186 11319 14188 11328
rect 14240 11319 14242 11328
rect 14188 11290 14240 11296
rect 14200 10810 14228 11290
rect 14188 10804 14240 10810
rect 14188 10746 14240 10752
rect 14188 10668 14240 10674
rect 14188 10610 14240 10616
rect 14200 10266 14228 10610
rect 14188 10260 14240 10266
rect 14188 10202 14240 10208
rect 14186 10160 14242 10169
rect 14186 10095 14242 10104
rect 14200 9897 14228 10095
rect 14186 9888 14242 9897
rect 14186 9823 14242 9832
rect 14200 9592 14228 9823
rect 14188 9586 14240 9592
rect 14188 9528 14240 9534
rect 14292 9500 14320 11999
rect 14384 11694 14412 14062
rect 14568 13802 14596 16623
rect 14556 13796 14608 13802
rect 14476 13756 14556 13784
rect 14372 11688 14424 11694
rect 14372 11630 14424 11636
rect 14384 11529 14412 11630
rect 14370 11520 14426 11529
rect 14370 11455 14426 11464
rect 14372 11144 14424 11150
rect 14372 11086 14424 11092
rect 14200 9472 14320 9500
rect 14200 9194 14228 9472
rect 14280 9376 14332 9382
rect 14278 9344 14280 9353
rect 14332 9344 14334 9353
rect 14278 9279 14334 9288
rect 14200 9166 14320 9194
rect 14188 8968 14240 8974
rect 14188 8910 14240 8916
rect 14096 6452 14148 6458
rect 14096 6394 14148 6400
rect 14200 6338 14228 8910
rect 14108 6310 14228 6338
rect 14004 5772 14056 5778
rect 14004 5714 14056 5720
rect 13912 4140 13964 4146
rect 13912 4082 13964 4088
rect 14016 3602 14044 5714
rect 14004 3596 14056 3602
rect 14004 3538 14056 3544
rect 14108 3194 14136 6310
rect 14186 5672 14242 5681
rect 14186 5607 14242 5616
rect 14200 5574 14228 5607
rect 14188 5568 14240 5574
rect 14188 5510 14240 5516
rect 14292 3992 14320 9166
rect 14384 7410 14412 11086
rect 14476 10606 14504 13756
rect 14556 13738 14608 13744
rect 14660 13410 14688 18294
rect 15292 18080 15344 18086
rect 15292 18022 15344 18028
rect 15200 16652 15252 16658
rect 15200 16594 15252 16600
rect 15212 16561 15240 16594
rect 15198 16552 15254 16561
rect 15198 16487 15254 16496
rect 14830 15736 14886 15745
rect 14830 15671 14886 15680
rect 14844 15638 14872 15671
rect 14832 15632 14884 15638
rect 14832 15574 14884 15580
rect 14740 14952 14792 14958
rect 14740 14894 14792 14900
rect 14752 13841 14780 14894
rect 14738 13832 14794 13841
rect 14738 13767 14794 13776
rect 14660 13382 14780 13410
rect 14648 13320 14700 13326
rect 14648 13262 14700 13268
rect 14660 12374 14688 13262
rect 14648 12368 14700 12374
rect 14554 12336 14610 12345
rect 14648 12310 14700 12316
rect 14554 12271 14610 12280
rect 14568 12186 14596 12271
rect 14568 12158 14688 12186
rect 14660 12102 14688 12158
rect 14556 12096 14608 12102
rect 14556 12038 14608 12044
rect 14648 12096 14700 12102
rect 14648 12038 14700 12044
rect 14568 10849 14596 12038
rect 14648 11688 14700 11694
rect 14648 11630 14700 11636
rect 14554 10840 14610 10849
rect 14554 10775 14610 10784
rect 14464 10600 14516 10606
rect 14464 10542 14516 10548
rect 14568 10538 14596 10775
rect 14556 10532 14608 10538
rect 14556 10474 14608 10480
rect 14462 10296 14518 10305
rect 14462 10231 14518 10240
rect 14476 9586 14504 10231
rect 14554 10160 14610 10169
rect 14554 10095 14610 10104
rect 14464 9580 14516 9586
rect 14464 9522 14516 9528
rect 14464 9444 14516 9450
rect 14464 9386 14516 9392
rect 14476 9353 14504 9386
rect 14462 9344 14518 9353
rect 14462 9279 14518 9288
rect 14464 9172 14516 9178
rect 14464 9114 14516 9120
rect 14476 7410 14504 9114
rect 14568 8537 14596 10095
rect 14554 8528 14610 8537
rect 14554 8463 14610 8472
rect 14556 8356 14608 8362
rect 14556 8298 14608 8304
rect 14372 7404 14424 7410
rect 14372 7346 14424 7352
rect 14464 7404 14516 7410
rect 14464 7346 14516 7352
rect 14384 7256 14412 7346
rect 14384 7228 14504 7256
rect 14370 7168 14426 7177
rect 14370 7103 14426 7112
rect 14384 4010 14412 7103
rect 14476 6118 14504 7228
rect 14464 6112 14516 6118
rect 14464 6054 14516 6060
rect 14464 5772 14516 5778
rect 14568 5760 14596 8298
rect 14660 6254 14688 11630
rect 14752 11354 14780 13382
rect 14844 12850 14872 15574
rect 15016 15496 15068 15502
rect 15016 15438 15068 15444
rect 14924 13728 14976 13734
rect 14924 13670 14976 13676
rect 14832 12844 14884 12850
rect 14832 12786 14884 12792
rect 14832 12436 14884 12442
rect 14832 12378 14884 12384
rect 14844 11626 14872 12378
rect 14832 11620 14884 11626
rect 14832 11562 14884 11568
rect 14844 11529 14872 11562
rect 14830 11520 14886 11529
rect 14830 11455 14886 11464
rect 14740 11348 14792 11354
rect 14740 11290 14792 11296
rect 14752 9586 14780 11290
rect 14830 10840 14886 10849
rect 14830 10775 14886 10784
rect 14844 10742 14872 10775
rect 14832 10736 14884 10742
rect 14832 10678 14884 10684
rect 14832 10600 14884 10606
rect 14832 10542 14884 10548
rect 14844 9926 14872 10542
rect 14832 9920 14884 9926
rect 14832 9862 14884 9868
rect 14740 9580 14792 9586
rect 14740 9522 14792 9528
rect 14740 9376 14792 9382
rect 14740 9318 14792 9324
rect 14752 7177 14780 9318
rect 14844 7970 14872 9862
rect 14936 9110 14964 13670
rect 15028 12986 15056 15438
rect 15200 15360 15252 15366
rect 15200 15302 15252 15308
rect 15108 14884 15160 14890
rect 15108 14826 15160 14832
rect 15016 12980 15068 12986
rect 15016 12922 15068 12928
rect 15016 12844 15068 12850
rect 15016 12786 15068 12792
rect 14924 9104 14976 9110
rect 14924 9046 14976 9052
rect 14922 8800 14978 8809
rect 14922 8735 14978 8744
rect 14936 8294 14964 8735
rect 14924 8288 14976 8294
rect 14924 8230 14976 8236
rect 14844 7942 14964 7970
rect 14832 7880 14884 7886
rect 14832 7822 14884 7828
rect 14844 7721 14872 7822
rect 14830 7712 14886 7721
rect 14830 7647 14886 7656
rect 14738 7168 14794 7177
rect 14738 7103 14794 7112
rect 14832 6928 14884 6934
rect 14832 6870 14884 6876
rect 14740 6656 14792 6662
rect 14740 6598 14792 6604
rect 14648 6248 14700 6254
rect 14648 6190 14700 6196
rect 14648 6112 14700 6118
rect 14648 6054 14700 6060
rect 14516 5732 14596 5760
rect 14464 5714 14516 5720
rect 14200 3964 14320 3992
rect 14372 4004 14424 4010
rect 14096 3188 14148 3194
rect 14096 3130 14148 3136
rect 14200 2854 14228 3964
rect 14372 3946 14424 3952
rect 14476 3890 14504 5714
rect 14554 5128 14610 5137
rect 14554 5063 14610 5072
rect 14568 4622 14596 5063
rect 14660 4826 14688 6054
rect 14648 4820 14700 4826
rect 14648 4762 14700 4768
rect 14646 4720 14702 4729
rect 14646 4655 14702 4664
rect 14660 4622 14688 4655
rect 14752 4622 14780 6598
rect 14844 5778 14872 6870
rect 14936 6186 14964 7942
rect 14924 6180 14976 6186
rect 14924 6122 14976 6128
rect 14832 5772 14884 5778
rect 14832 5714 14884 5720
rect 14924 5636 14976 5642
rect 14924 5578 14976 5584
rect 14832 5568 14884 5574
rect 14832 5510 14884 5516
rect 14844 4865 14872 5510
rect 14830 4856 14886 4865
rect 14830 4791 14886 4800
rect 14844 4758 14872 4791
rect 14832 4752 14884 4758
rect 14832 4694 14884 4700
rect 14556 4616 14608 4622
rect 14556 4558 14608 4564
rect 14648 4616 14700 4622
rect 14648 4558 14700 4564
rect 14740 4616 14792 4622
rect 14740 4558 14792 4564
rect 14292 3862 14504 3890
rect 14292 3176 14320 3862
rect 14464 3188 14516 3194
rect 14292 3148 14464 3176
rect 14188 2848 14240 2854
rect 14188 2790 14240 2796
rect 13820 2508 13872 2514
rect 13820 2450 13872 2456
rect 13728 2440 13780 2446
rect 13728 2382 13780 2388
rect 13544 2032 13596 2038
rect 13544 1974 13596 1980
rect 13084 1488 13136 1494
rect 13084 1430 13136 1436
rect 12992 1284 13044 1290
rect 12992 1226 13044 1232
rect 12532 672 12584 678
rect 11610 640 11666 649
rect 12532 614 12584 620
rect 14292 610 14320 3148
rect 14464 3130 14516 3136
rect 11610 575 11666 584
rect 14280 604 14332 610
rect 14280 546 14332 552
rect 14660 542 14688 4558
rect 14936 4146 14964 5578
rect 15028 4622 15056 12786
rect 15120 12442 15148 14826
rect 15212 14822 15240 15302
rect 15200 14816 15252 14822
rect 15200 14758 15252 14764
rect 15200 13320 15252 13326
rect 15200 13262 15252 13268
rect 15108 12436 15160 12442
rect 15108 12378 15160 12384
rect 15108 11008 15160 11014
rect 15108 10950 15160 10956
rect 15120 10810 15148 10950
rect 15108 10804 15160 10810
rect 15108 10746 15160 10752
rect 15212 10724 15240 13262
rect 15304 12986 15332 18022
rect 15948 17814 15976 18498
rect 15936 17808 15988 17814
rect 15936 17750 15988 17756
rect 15384 17604 15436 17610
rect 15384 17546 15436 17552
rect 15292 12980 15344 12986
rect 15292 12922 15344 12928
rect 15396 12238 15424 17546
rect 15660 17332 15712 17338
rect 15660 17274 15712 17280
rect 15568 16788 15620 16794
rect 15568 16730 15620 16736
rect 15476 13320 15528 13326
rect 15474 13288 15476 13297
rect 15528 13288 15530 13297
rect 15474 13223 15530 13232
rect 15476 12980 15528 12986
rect 15476 12922 15528 12928
rect 15384 12232 15436 12238
rect 15384 12174 15436 12180
rect 15292 12164 15344 12170
rect 15292 12106 15344 12112
rect 15304 10849 15332 12106
rect 15290 10840 15346 10849
rect 15290 10775 15346 10784
rect 15212 10696 15332 10724
rect 15108 10668 15160 10674
rect 15108 10610 15160 10616
rect 15120 10198 15148 10610
rect 15198 10296 15254 10305
rect 15198 10231 15254 10240
rect 15108 10192 15160 10198
rect 15108 10134 15160 10140
rect 15108 10056 15160 10062
rect 15108 9998 15160 10004
rect 15120 9722 15148 9998
rect 15108 9716 15160 9722
rect 15108 9658 15160 9664
rect 15212 9674 15240 10231
rect 15304 10062 15332 10696
rect 15396 10470 15424 12174
rect 15488 11830 15516 12922
rect 15476 11824 15528 11830
rect 15476 11766 15528 11772
rect 15580 11014 15608 16730
rect 15672 12617 15700 17274
rect 16132 17202 16160 19200
rect 17498 18592 17554 18601
rect 17498 18527 17554 18536
rect 17406 18456 17462 18465
rect 16764 18420 16816 18426
rect 17406 18391 17462 18400
rect 16764 18362 16816 18368
rect 16304 18216 16356 18222
rect 16304 18158 16356 18164
rect 16120 17196 16172 17202
rect 16120 17138 16172 17144
rect 16028 17128 16080 17134
rect 16028 17070 16080 17076
rect 16040 14958 16068 17070
rect 16212 16720 16264 16726
rect 16212 16662 16264 16668
rect 16120 16584 16172 16590
rect 16120 16526 16172 16532
rect 16028 14952 16080 14958
rect 16028 14894 16080 14900
rect 15752 14612 15804 14618
rect 15752 14554 15804 14560
rect 15764 13938 15792 14554
rect 15936 14476 15988 14482
rect 15936 14418 15988 14424
rect 15752 13932 15804 13938
rect 15752 13874 15804 13880
rect 15658 12608 15714 12617
rect 15658 12543 15714 12552
rect 15764 12434 15792 13874
rect 15844 13184 15896 13190
rect 15844 13126 15896 13132
rect 15672 12406 15792 12434
rect 15672 11150 15700 12406
rect 15752 12368 15804 12374
rect 15752 12310 15804 12316
rect 15660 11144 15712 11150
rect 15660 11086 15712 11092
rect 15568 11008 15620 11014
rect 15568 10950 15620 10956
rect 15476 10804 15528 10810
rect 15476 10746 15528 10752
rect 15660 10804 15712 10810
rect 15660 10746 15712 10752
rect 15384 10464 15436 10470
rect 15384 10406 15436 10412
rect 15384 10260 15436 10266
rect 15384 10202 15436 10208
rect 15292 10056 15344 10062
rect 15292 9998 15344 10004
rect 15396 9994 15424 10202
rect 15384 9988 15436 9994
rect 15384 9930 15436 9936
rect 15488 9674 15516 10746
rect 15568 10668 15620 10674
rect 15568 10610 15620 10616
rect 15212 9646 15332 9674
rect 15106 9616 15162 9625
rect 15106 9551 15108 9560
rect 15160 9551 15162 9560
rect 15108 9522 15160 9528
rect 15200 9104 15252 9110
rect 15200 9046 15252 9052
rect 15108 8832 15160 8838
rect 15108 8774 15160 8780
rect 15120 8634 15148 8774
rect 15108 8628 15160 8634
rect 15108 8570 15160 8576
rect 15106 8120 15162 8129
rect 15106 8055 15162 8064
rect 15120 8022 15148 8055
rect 15108 8016 15160 8022
rect 15108 7958 15160 7964
rect 15120 7478 15148 7958
rect 15108 7472 15160 7478
rect 15108 7414 15160 7420
rect 15120 5846 15148 7414
rect 15108 5840 15160 5846
rect 15108 5782 15160 5788
rect 15212 5710 15240 9046
rect 15108 5704 15160 5710
rect 15108 5646 15160 5652
rect 15200 5704 15252 5710
rect 15200 5646 15252 5652
rect 15016 4616 15068 4622
rect 15016 4558 15068 4564
rect 14924 4140 14976 4146
rect 14924 4082 14976 4088
rect 15120 4010 15148 5646
rect 15200 5568 15252 5574
rect 15200 5510 15252 5516
rect 15212 4282 15240 5510
rect 15304 4826 15332 9646
rect 15396 9646 15516 9674
rect 15396 8616 15424 9646
rect 15476 9512 15528 9518
rect 15580 9489 15608 10610
rect 15476 9454 15528 9460
rect 15566 9480 15622 9489
rect 15488 9364 15516 9454
rect 15566 9415 15622 9424
rect 15488 9336 15608 9364
rect 15396 8588 15516 8616
rect 15384 8492 15436 8498
rect 15384 8434 15436 8440
rect 15396 7886 15424 8434
rect 15488 8430 15516 8588
rect 15476 8424 15528 8430
rect 15476 8366 15528 8372
rect 15476 8288 15528 8294
rect 15476 8230 15528 8236
rect 15488 7886 15516 8230
rect 15384 7880 15436 7886
rect 15384 7822 15436 7828
rect 15476 7880 15528 7886
rect 15476 7822 15528 7828
rect 15382 7032 15438 7041
rect 15382 6967 15438 6976
rect 15396 6769 15424 6967
rect 15382 6760 15438 6769
rect 15382 6695 15438 6704
rect 15292 4820 15344 4826
rect 15292 4762 15344 4768
rect 15200 4276 15252 4282
rect 15200 4218 15252 4224
rect 14924 4004 14976 4010
rect 14924 3946 14976 3952
rect 15108 4004 15160 4010
rect 15108 3946 15160 3952
rect 14936 1766 14964 3946
rect 15396 3942 15424 6695
rect 15488 6390 15516 7822
rect 15476 6384 15528 6390
rect 15476 6326 15528 6332
rect 15476 5228 15528 5234
rect 15476 5170 15528 5176
rect 15384 3936 15436 3942
rect 15384 3878 15436 3884
rect 15292 3596 15344 3602
rect 15292 3538 15344 3544
rect 15304 2632 15332 3538
rect 15384 3460 15436 3466
rect 15384 3402 15436 3408
rect 15396 3097 15424 3402
rect 15382 3088 15438 3097
rect 15382 3023 15438 3032
rect 15304 2604 15424 2632
rect 15292 2508 15344 2514
rect 15292 2450 15344 2456
rect 14924 1760 14976 1766
rect 14924 1702 14976 1708
rect 15304 1057 15332 2450
rect 15290 1048 15346 1057
rect 15290 983 15346 992
rect 15396 950 15424 2604
rect 15384 944 15436 950
rect 15384 886 15436 892
rect 15488 882 15516 5170
rect 15580 2961 15608 9336
rect 15672 8945 15700 10746
rect 15658 8936 15714 8945
rect 15658 8871 15714 8880
rect 15764 8566 15792 12310
rect 15856 11558 15884 13126
rect 15948 12782 15976 14418
rect 16040 14074 16068 14894
rect 16028 14068 16080 14074
rect 16028 14010 16080 14016
rect 16028 12980 16080 12986
rect 16028 12922 16080 12928
rect 16040 12850 16068 12922
rect 16028 12844 16080 12850
rect 16028 12786 16080 12792
rect 15936 12776 15988 12782
rect 15936 12718 15988 12724
rect 15934 12608 15990 12617
rect 15934 12543 15990 12552
rect 15948 12170 15976 12543
rect 15936 12164 15988 12170
rect 15936 12106 15988 12112
rect 16132 11812 16160 16526
rect 16224 12442 16252 16662
rect 16316 14278 16344 18158
rect 16488 17672 16540 17678
rect 16488 17614 16540 17620
rect 16396 16516 16448 16522
rect 16396 16458 16448 16464
rect 16408 15706 16436 16458
rect 16396 15700 16448 15706
rect 16396 15642 16448 15648
rect 16394 15056 16450 15065
rect 16394 14991 16450 15000
rect 16408 14414 16436 14991
rect 16500 14618 16528 17614
rect 16672 17536 16724 17542
rect 16672 17478 16724 17484
rect 16580 16108 16632 16114
rect 16580 16050 16632 16056
rect 16592 14906 16620 16050
rect 16684 15026 16712 17478
rect 16776 16538 16804 18362
rect 17314 17232 17370 17241
rect 17314 17167 17316 17176
rect 17368 17167 17370 17176
rect 17316 17138 17368 17144
rect 17316 17060 17368 17066
rect 17316 17002 17368 17008
rect 16950 16892 17258 16901
rect 16950 16890 16956 16892
rect 17012 16890 17036 16892
rect 17092 16890 17116 16892
rect 17172 16890 17196 16892
rect 17252 16890 17258 16892
rect 17012 16838 17014 16890
rect 17194 16838 17196 16890
rect 16950 16836 16956 16838
rect 17012 16836 17036 16838
rect 17092 16836 17116 16838
rect 17172 16836 17196 16838
rect 17252 16836 17258 16838
rect 16950 16827 17258 16836
rect 17040 16584 17092 16590
rect 16776 16510 16896 16538
rect 17132 16584 17184 16590
rect 17040 16526 17092 16532
rect 17130 16552 17132 16561
rect 17184 16552 17186 16561
rect 16764 16448 16816 16454
rect 16764 16390 16816 16396
rect 16776 15570 16804 16390
rect 16764 15564 16816 15570
rect 16764 15506 16816 15512
rect 16672 15020 16724 15026
rect 16672 14962 16724 14968
rect 16592 14878 16804 14906
rect 16488 14612 16540 14618
rect 16488 14554 16540 14560
rect 16500 14482 16528 14554
rect 16488 14476 16540 14482
rect 16488 14418 16540 14424
rect 16396 14408 16448 14414
rect 16672 14408 16724 14414
rect 16396 14350 16448 14356
rect 16592 14368 16672 14396
rect 16304 14272 16356 14278
rect 16304 14214 16356 14220
rect 16302 13016 16358 13025
rect 16302 12951 16358 12960
rect 16316 12918 16344 12951
rect 16304 12912 16356 12918
rect 16304 12854 16356 12860
rect 16408 12458 16436 14350
rect 16592 13870 16620 14368
rect 16672 14350 16724 14356
rect 16776 14278 16804 14878
rect 16672 14272 16724 14278
rect 16672 14214 16724 14220
rect 16764 14272 16816 14278
rect 16764 14214 16816 14220
rect 16580 13864 16632 13870
rect 16580 13806 16632 13812
rect 16684 13326 16712 14214
rect 16868 13512 16896 16510
rect 17052 16153 17080 16526
rect 17130 16487 17186 16496
rect 17144 16250 17172 16487
rect 17132 16244 17184 16250
rect 17132 16186 17184 16192
rect 17038 16144 17094 16153
rect 17038 16079 17094 16088
rect 16950 15804 17258 15813
rect 16950 15802 16956 15804
rect 17012 15802 17036 15804
rect 17092 15802 17116 15804
rect 17172 15802 17196 15804
rect 17252 15802 17258 15804
rect 17012 15750 17014 15802
rect 17194 15750 17196 15802
rect 16950 15748 16956 15750
rect 17012 15748 17036 15750
rect 17092 15748 17116 15750
rect 17172 15748 17196 15750
rect 17252 15748 17258 15750
rect 16950 15739 17258 15748
rect 16950 14716 17258 14725
rect 16950 14714 16956 14716
rect 17012 14714 17036 14716
rect 17092 14714 17116 14716
rect 17172 14714 17196 14716
rect 17252 14714 17258 14716
rect 17012 14662 17014 14714
rect 17194 14662 17196 14714
rect 16950 14660 16956 14662
rect 17012 14660 17036 14662
rect 17092 14660 17116 14662
rect 17172 14660 17196 14662
rect 17252 14660 17258 14662
rect 16950 14651 17258 14660
rect 17132 14272 17184 14278
rect 17132 14214 17184 14220
rect 17144 13734 17172 14214
rect 17132 13728 17184 13734
rect 17132 13670 17184 13676
rect 16950 13628 17258 13637
rect 16950 13626 16956 13628
rect 17012 13626 17036 13628
rect 17092 13626 17116 13628
rect 17172 13626 17196 13628
rect 17252 13626 17258 13628
rect 17012 13574 17014 13626
rect 17194 13574 17196 13626
rect 16950 13572 16956 13574
rect 17012 13572 17036 13574
rect 17092 13572 17116 13574
rect 17172 13572 17196 13574
rect 17252 13572 17258 13574
rect 16950 13563 17258 13572
rect 17224 13524 17276 13530
rect 16868 13484 16988 13512
rect 16672 13320 16724 13326
rect 16672 13262 16724 13268
rect 16856 13252 16908 13258
rect 16856 13194 16908 13200
rect 16868 12696 16896 13194
rect 16776 12668 16896 12696
rect 16212 12436 16264 12442
rect 16408 12430 16620 12458
rect 16212 12378 16264 12384
rect 16488 12368 16540 12374
rect 16408 12328 16488 12356
rect 16304 12232 16356 12238
rect 16304 12174 16356 12180
rect 16040 11784 16160 11812
rect 15936 11688 15988 11694
rect 15936 11630 15988 11636
rect 15844 11552 15896 11558
rect 15844 11494 15896 11500
rect 15844 11280 15896 11286
rect 15842 11248 15844 11257
rect 15896 11248 15898 11257
rect 15842 11183 15898 11192
rect 15856 11150 15884 11183
rect 15844 11144 15896 11150
rect 15844 11086 15896 11092
rect 15948 10849 15976 11630
rect 15934 10840 15990 10849
rect 15934 10775 15990 10784
rect 15844 10464 15896 10470
rect 15844 10406 15896 10412
rect 15934 10432 15990 10441
rect 15856 10305 15884 10406
rect 15934 10367 15990 10376
rect 15842 10296 15898 10305
rect 15842 10231 15898 10240
rect 15844 10192 15896 10198
rect 15844 10134 15896 10140
rect 15752 8560 15804 8566
rect 15752 8502 15804 8508
rect 15660 8424 15712 8430
rect 15660 8366 15712 8372
rect 15672 6338 15700 8366
rect 15856 8106 15884 10134
rect 15948 9586 15976 10367
rect 15936 9580 15988 9586
rect 15936 9522 15988 9528
rect 15936 9444 15988 9450
rect 15936 9386 15988 9392
rect 15764 8078 15884 8106
rect 15764 7342 15792 8078
rect 15844 8016 15896 8022
rect 15844 7958 15896 7964
rect 15856 7750 15884 7958
rect 15844 7744 15896 7750
rect 15844 7686 15896 7692
rect 15752 7336 15804 7342
rect 15752 7278 15804 7284
rect 15856 7002 15884 7686
rect 15844 6996 15896 7002
rect 15844 6938 15896 6944
rect 15948 6458 15976 9386
rect 16040 8090 16068 11784
rect 16212 10668 16264 10674
rect 16132 10628 16212 10656
rect 16132 10266 16160 10628
rect 16212 10610 16264 10616
rect 16316 10554 16344 12174
rect 16224 10526 16344 10554
rect 16120 10260 16172 10266
rect 16120 10202 16172 10208
rect 16224 9976 16252 10526
rect 16304 10464 16356 10470
rect 16304 10406 16356 10412
rect 16316 10112 16344 10406
rect 16132 9948 16252 9976
rect 16292 10084 16344 10112
rect 16028 8084 16080 8090
rect 16028 8026 16080 8032
rect 16132 7970 16160 9948
rect 16292 9874 16320 10084
rect 16292 9846 16344 9874
rect 16212 9512 16264 9518
rect 16316 9500 16344 9846
rect 16264 9472 16344 9500
rect 16212 9454 16264 9460
rect 16304 9376 16356 9382
rect 16304 9318 16356 9324
rect 16040 7942 16160 7970
rect 16210 7984 16266 7993
rect 15936 6452 15988 6458
rect 15936 6394 15988 6400
rect 16040 6361 16068 7942
rect 16210 7919 16212 7928
rect 16264 7919 16266 7928
rect 16212 7890 16264 7896
rect 16120 7880 16172 7886
rect 16316 7834 16344 9318
rect 16408 9042 16436 12328
rect 16488 12310 16540 12316
rect 16488 12232 16540 12238
rect 16486 12200 16488 12209
rect 16592 12220 16620 12430
rect 16672 12232 16724 12238
rect 16540 12200 16542 12209
rect 16592 12192 16672 12220
rect 16672 12174 16724 12180
rect 16486 12135 16542 12144
rect 16488 11892 16540 11898
rect 16488 11834 16540 11840
rect 16500 11082 16528 11834
rect 16580 11824 16632 11830
rect 16580 11766 16632 11772
rect 16670 11792 16726 11801
rect 16488 11076 16540 11082
rect 16488 11018 16540 11024
rect 16500 10266 16528 11018
rect 16488 10260 16540 10266
rect 16488 10202 16540 10208
rect 16488 10056 16540 10062
rect 16488 9998 16540 10004
rect 16500 9761 16528 9998
rect 16486 9752 16542 9761
rect 16486 9687 16542 9696
rect 16592 9674 16620 11766
rect 16670 11727 16726 11736
rect 16684 9994 16712 11727
rect 16776 11694 16804 12668
rect 16960 12628 16988 13484
rect 17224 13466 17276 13472
rect 17236 12850 17264 13466
rect 17224 12844 17276 12850
rect 17224 12786 17276 12792
rect 16868 12600 16988 12628
rect 16868 11830 16896 12600
rect 16950 12540 17258 12549
rect 16950 12538 16956 12540
rect 17012 12538 17036 12540
rect 17092 12538 17116 12540
rect 17172 12538 17196 12540
rect 17252 12538 17258 12540
rect 17012 12486 17014 12538
rect 17194 12486 17196 12538
rect 16950 12484 16956 12486
rect 17012 12484 17036 12486
rect 17092 12484 17116 12486
rect 17172 12484 17196 12486
rect 17252 12484 17258 12486
rect 16950 12475 17258 12484
rect 16948 12300 17000 12306
rect 16948 12242 17000 12248
rect 16856 11824 16908 11830
rect 16856 11766 16908 11772
rect 16764 11688 16816 11694
rect 16960 11676 16988 12242
rect 17040 12232 17092 12238
rect 17040 12174 17092 12180
rect 17052 11898 17080 12174
rect 17040 11892 17092 11898
rect 17040 11834 17092 11840
rect 16764 11630 16816 11636
rect 16868 11648 16988 11676
rect 16764 11552 16816 11558
rect 16764 11494 16816 11500
rect 16776 10266 16804 11494
rect 16868 11218 16896 11648
rect 16950 11452 17258 11461
rect 16950 11450 16956 11452
rect 17012 11450 17036 11452
rect 17092 11450 17116 11452
rect 17172 11450 17196 11452
rect 17252 11450 17258 11452
rect 17012 11398 17014 11450
rect 17194 11398 17196 11450
rect 16950 11396 16956 11398
rect 17012 11396 17036 11398
rect 17092 11396 17116 11398
rect 17172 11396 17196 11398
rect 17252 11396 17258 11398
rect 16950 11387 17258 11396
rect 16948 11348 17000 11354
rect 16948 11290 17000 11296
rect 16856 11212 16908 11218
rect 16856 11154 16908 11160
rect 16960 10742 16988 11290
rect 17038 10976 17094 10985
rect 17038 10911 17094 10920
rect 16948 10736 17000 10742
rect 16948 10678 17000 10684
rect 17052 10606 17080 10911
rect 17040 10600 17092 10606
rect 17040 10542 17092 10548
rect 17040 10464 17092 10470
rect 16868 10424 17040 10452
rect 16764 10260 16816 10266
rect 16764 10202 16816 10208
rect 16762 10160 16818 10169
rect 16762 10095 16818 10104
rect 16672 9988 16724 9994
rect 16672 9930 16724 9936
rect 16592 9646 16712 9674
rect 16486 9616 16542 9625
rect 16486 9551 16488 9560
rect 16540 9551 16542 9560
rect 16488 9522 16540 9528
rect 16684 9466 16712 9646
rect 16488 9444 16540 9450
rect 16488 9386 16540 9392
rect 16592 9438 16712 9466
rect 16396 9036 16448 9042
rect 16396 8978 16448 8984
rect 16500 8906 16528 9386
rect 16488 8900 16540 8906
rect 16488 8842 16540 8848
rect 16396 8832 16448 8838
rect 16448 8780 16528 8786
rect 16396 8774 16528 8780
rect 16408 8758 16528 8774
rect 16396 8628 16448 8634
rect 16396 8570 16448 8576
rect 16120 7822 16172 7828
rect 16026 6352 16082 6361
rect 15672 6310 15884 6338
rect 15752 6180 15804 6186
rect 15752 6122 15804 6128
rect 15660 5228 15712 5234
rect 15660 5170 15712 5176
rect 15672 4185 15700 5170
rect 15658 4176 15714 4185
rect 15658 4111 15714 4120
rect 15764 3602 15792 6122
rect 15752 3596 15804 3602
rect 15752 3538 15804 3544
rect 15856 3482 15884 6310
rect 16026 6287 16082 6296
rect 16028 5840 16080 5846
rect 16028 5782 16080 5788
rect 15934 5536 15990 5545
rect 15934 5471 15990 5480
rect 15948 4690 15976 5471
rect 15936 4684 15988 4690
rect 15936 4626 15988 4632
rect 15948 4457 15976 4626
rect 15934 4448 15990 4457
rect 15934 4383 15990 4392
rect 16040 4298 16068 5782
rect 16132 5166 16160 7822
rect 16224 7806 16344 7834
rect 16224 6633 16252 7806
rect 16304 7744 16356 7750
rect 16304 7686 16356 7692
rect 16316 7546 16344 7686
rect 16304 7540 16356 7546
rect 16304 7482 16356 7488
rect 16210 6624 16266 6633
rect 16210 6559 16266 6568
rect 16210 6488 16266 6497
rect 16210 6423 16266 6432
rect 16120 5160 16172 5166
rect 16120 5102 16172 5108
rect 16120 4616 16172 4622
rect 16120 4558 16172 4564
rect 15948 4270 16068 4298
rect 15948 3602 15976 4270
rect 16026 4176 16082 4185
rect 16026 4111 16082 4120
rect 15936 3596 15988 3602
rect 15936 3538 15988 3544
rect 16040 3534 16068 4111
rect 15672 3454 15884 3482
rect 16028 3528 16080 3534
rect 16028 3470 16080 3476
rect 15566 2952 15622 2961
rect 15566 2887 15622 2896
rect 15672 2378 15700 3454
rect 15844 3052 15896 3058
rect 15844 2994 15896 3000
rect 15660 2372 15712 2378
rect 15660 2314 15712 2320
rect 15856 921 15884 2994
rect 16040 1086 16068 3470
rect 16132 3369 16160 4558
rect 16118 3360 16174 3369
rect 16118 3295 16174 3304
rect 16224 3126 16252 6423
rect 16304 5704 16356 5710
rect 16304 5646 16356 5652
rect 16316 4622 16344 5646
rect 16408 5370 16436 8570
rect 16500 6089 16528 8758
rect 16592 6118 16620 9438
rect 16776 9110 16804 10095
rect 16764 9104 16816 9110
rect 16764 9046 16816 9052
rect 16672 8968 16724 8974
rect 16672 8910 16724 8916
rect 16580 6112 16632 6118
rect 16486 6080 16542 6089
rect 16580 6054 16632 6060
rect 16486 6015 16542 6024
rect 16578 5944 16634 5953
rect 16578 5879 16634 5888
rect 16592 5778 16620 5879
rect 16488 5772 16540 5778
rect 16488 5714 16540 5720
rect 16580 5772 16632 5778
rect 16580 5714 16632 5720
rect 16396 5364 16448 5370
rect 16396 5306 16448 5312
rect 16500 5302 16528 5714
rect 16580 5636 16632 5642
rect 16580 5578 16632 5584
rect 16488 5296 16540 5302
rect 16488 5238 16540 5244
rect 16488 5160 16540 5166
rect 16488 5102 16540 5108
rect 16304 4616 16356 4622
rect 16304 4558 16356 4564
rect 16302 4448 16358 4457
rect 16302 4383 16358 4392
rect 16316 3466 16344 4383
rect 16396 4208 16448 4214
rect 16396 4150 16448 4156
rect 16408 3738 16436 4150
rect 16396 3732 16448 3738
rect 16396 3674 16448 3680
rect 16408 3534 16436 3674
rect 16396 3528 16448 3534
rect 16396 3470 16448 3476
rect 16304 3460 16356 3466
rect 16304 3402 16356 3408
rect 16212 3120 16264 3126
rect 16212 3062 16264 3068
rect 16500 3058 16528 5102
rect 16592 3738 16620 5578
rect 16684 5166 16712 8910
rect 16764 8832 16816 8838
rect 16764 8774 16816 8780
rect 16776 8090 16804 8774
rect 16764 8084 16816 8090
rect 16764 8026 16816 8032
rect 16868 6916 16896 10424
rect 17040 10406 17092 10412
rect 16950 10364 17258 10373
rect 16950 10362 16956 10364
rect 17012 10362 17036 10364
rect 17092 10362 17116 10364
rect 17172 10362 17196 10364
rect 17252 10362 17258 10364
rect 17012 10310 17014 10362
rect 17194 10310 17196 10362
rect 16950 10308 16956 10310
rect 17012 10308 17036 10310
rect 17092 10308 17116 10310
rect 17172 10308 17196 10310
rect 17252 10308 17258 10310
rect 16950 10299 17258 10308
rect 16948 10260 17000 10266
rect 16948 10202 17000 10208
rect 16960 9654 16988 10202
rect 17040 10056 17092 10062
rect 17040 9998 17092 10004
rect 17052 9897 17080 9998
rect 17038 9888 17094 9897
rect 17038 9823 17094 9832
rect 17224 9716 17276 9722
rect 17224 9658 17276 9664
rect 16948 9648 17000 9654
rect 16948 9590 17000 9596
rect 17236 9586 17264 9658
rect 17224 9580 17276 9586
rect 17224 9522 17276 9528
rect 16950 9276 17258 9285
rect 16950 9274 16956 9276
rect 17012 9274 17036 9276
rect 17092 9274 17116 9276
rect 17172 9274 17196 9276
rect 17252 9274 17258 9276
rect 17012 9222 17014 9274
rect 17194 9222 17196 9274
rect 16950 9220 16956 9222
rect 17012 9220 17036 9222
rect 17092 9220 17116 9222
rect 17172 9220 17196 9222
rect 17252 9220 17258 9222
rect 16950 9211 17258 9220
rect 17224 9104 17276 9110
rect 17224 9046 17276 9052
rect 17236 8974 17264 9046
rect 17224 8968 17276 8974
rect 17224 8910 17276 8916
rect 16950 8188 17258 8197
rect 16950 8186 16956 8188
rect 17012 8186 17036 8188
rect 17092 8186 17116 8188
rect 17172 8186 17196 8188
rect 17252 8186 17258 8188
rect 17012 8134 17014 8186
rect 17194 8134 17196 8186
rect 16950 8132 16956 8134
rect 17012 8132 17036 8134
rect 17092 8132 17116 8134
rect 17172 8132 17196 8134
rect 17252 8132 17258 8134
rect 16950 8123 17258 8132
rect 17040 7880 17092 7886
rect 17038 7848 17040 7857
rect 17092 7848 17094 7857
rect 17038 7783 17094 7792
rect 17224 7812 17276 7818
rect 17224 7754 17276 7760
rect 17236 7478 17264 7754
rect 17224 7472 17276 7478
rect 17224 7414 17276 7420
rect 17040 7404 17092 7410
rect 17040 7346 17092 7352
rect 17052 7313 17080 7346
rect 17038 7304 17094 7313
rect 17038 7239 17094 7248
rect 16950 7100 17258 7109
rect 16950 7098 16956 7100
rect 17012 7098 17036 7100
rect 17092 7098 17116 7100
rect 17172 7098 17196 7100
rect 17252 7098 17258 7100
rect 17012 7046 17014 7098
rect 17194 7046 17196 7098
rect 16950 7044 16956 7046
rect 17012 7044 17036 7046
rect 17092 7044 17116 7046
rect 17172 7044 17196 7046
rect 17252 7044 17258 7046
rect 16950 7035 17258 7044
rect 16776 6888 16896 6916
rect 16776 6225 16804 6888
rect 16856 6724 16908 6730
rect 16856 6666 16908 6672
rect 16762 6216 16818 6225
rect 16762 6151 16818 6160
rect 16868 5914 16896 6666
rect 16950 6012 17258 6021
rect 16950 6010 16956 6012
rect 17012 6010 17036 6012
rect 17092 6010 17116 6012
rect 17172 6010 17196 6012
rect 17252 6010 17258 6012
rect 17012 5958 17014 6010
rect 17194 5958 17196 6010
rect 16950 5956 16956 5958
rect 17012 5956 17036 5958
rect 17092 5956 17116 5958
rect 17172 5956 17196 5958
rect 17252 5956 17258 5958
rect 16950 5947 17258 5956
rect 16856 5908 16908 5914
rect 16856 5850 16908 5856
rect 17328 5778 17356 17002
rect 17420 15026 17448 18391
rect 17512 17338 17540 18527
rect 18326 17776 18382 17785
rect 18326 17711 18382 17720
rect 17610 17436 17918 17445
rect 17610 17434 17616 17436
rect 17672 17434 17696 17436
rect 17752 17434 17776 17436
rect 17832 17434 17856 17436
rect 17912 17434 17918 17436
rect 17672 17382 17674 17434
rect 17854 17382 17856 17434
rect 17610 17380 17616 17382
rect 17672 17380 17696 17382
rect 17752 17380 17776 17382
rect 17832 17380 17856 17382
rect 17912 17380 17918 17382
rect 17610 17371 17918 17380
rect 17500 17332 17552 17338
rect 17500 17274 17552 17280
rect 18144 17128 18196 17134
rect 18144 17070 18196 17076
rect 17960 16516 18012 16522
rect 17960 16458 18012 16464
rect 17610 16348 17918 16357
rect 17610 16346 17616 16348
rect 17672 16346 17696 16348
rect 17752 16346 17776 16348
rect 17832 16346 17856 16348
rect 17912 16346 17918 16348
rect 17672 16294 17674 16346
rect 17854 16294 17856 16346
rect 17610 16292 17616 16294
rect 17672 16292 17696 16294
rect 17752 16292 17776 16294
rect 17832 16292 17856 16294
rect 17912 16292 17918 16294
rect 17610 16283 17918 16292
rect 17500 16040 17552 16046
rect 17500 15982 17552 15988
rect 17408 15020 17460 15026
rect 17408 14962 17460 14968
rect 17512 14906 17540 15982
rect 17610 15260 17918 15269
rect 17610 15258 17616 15260
rect 17672 15258 17696 15260
rect 17752 15258 17776 15260
rect 17832 15258 17856 15260
rect 17912 15258 17918 15260
rect 17672 15206 17674 15258
rect 17854 15206 17856 15258
rect 17610 15204 17616 15206
rect 17672 15204 17696 15206
rect 17752 15204 17776 15206
rect 17832 15204 17856 15206
rect 17912 15204 17918 15206
rect 17610 15195 17918 15204
rect 17420 14878 17540 14906
rect 17420 12646 17448 14878
rect 17500 14544 17552 14550
rect 17500 14486 17552 14492
rect 17512 13569 17540 14486
rect 17610 14172 17918 14181
rect 17610 14170 17616 14172
rect 17672 14170 17696 14172
rect 17752 14170 17776 14172
rect 17832 14170 17856 14172
rect 17912 14170 17918 14172
rect 17672 14118 17674 14170
rect 17854 14118 17856 14170
rect 17610 14116 17616 14118
rect 17672 14116 17696 14118
rect 17752 14116 17776 14118
rect 17832 14116 17856 14118
rect 17912 14116 17918 14118
rect 17610 14107 17918 14116
rect 17498 13560 17554 13569
rect 17498 13495 17554 13504
rect 17500 13252 17552 13258
rect 17500 13194 17552 13200
rect 17408 12640 17460 12646
rect 17408 12582 17460 12588
rect 17512 12442 17540 13194
rect 17610 13084 17918 13093
rect 17610 13082 17616 13084
rect 17672 13082 17696 13084
rect 17752 13082 17776 13084
rect 17832 13082 17856 13084
rect 17912 13082 17918 13084
rect 17672 13030 17674 13082
rect 17854 13030 17856 13082
rect 17610 13028 17616 13030
rect 17672 13028 17696 13030
rect 17752 13028 17776 13030
rect 17832 13028 17856 13030
rect 17912 13028 17918 13030
rect 17610 13019 17918 13028
rect 17682 12880 17738 12889
rect 17682 12815 17684 12824
rect 17736 12815 17738 12824
rect 17684 12786 17736 12792
rect 17682 12744 17738 12753
rect 17682 12679 17738 12688
rect 17500 12436 17552 12442
rect 17500 12378 17552 12384
rect 17408 12300 17460 12306
rect 17460 12260 17540 12288
rect 17408 12242 17460 12248
rect 17406 11928 17462 11937
rect 17406 11863 17462 11872
rect 17420 11762 17448 11863
rect 17408 11756 17460 11762
rect 17408 11698 17460 11704
rect 17512 11642 17540 12260
rect 17696 12186 17724 12679
rect 17972 12288 18000 16458
rect 18156 15609 18184 17070
rect 18236 16176 18288 16182
rect 18236 16118 18288 16124
rect 18142 15600 18198 15609
rect 18142 15535 18198 15544
rect 18156 15026 18184 15535
rect 18144 15020 18196 15026
rect 18144 14962 18196 14968
rect 18248 14906 18276 16118
rect 18156 14878 18276 14906
rect 18052 14340 18104 14346
rect 18052 14282 18104 14288
rect 18064 12986 18092 14282
rect 18052 12980 18104 12986
rect 18052 12922 18104 12928
rect 18156 12374 18184 14878
rect 18236 14408 18288 14414
rect 18236 14350 18288 14356
rect 18248 13938 18276 14350
rect 18236 13932 18288 13938
rect 18236 13874 18288 13880
rect 18236 13320 18288 13326
rect 18236 13262 18288 13268
rect 18248 12889 18276 13262
rect 18340 12918 18368 17711
rect 18616 17202 18644 19200
rect 19524 17808 19576 17814
rect 19524 17750 19576 17756
rect 18604 17196 18656 17202
rect 18604 17138 18656 17144
rect 18420 16448 18472 16454
rect 18420 16390 18472 16396
rect 18432 16153 18460 16390
rect 18418 16144 18474 16153
rect 18418 16079 18474 16088
rect 18788 15904 18840 15910
rect 18788 15846 18840 15852
rect 18418 13696 18474 13705
rect 18418 13631 18474 13640
rect 18432 13530 18460 13631
rect 18420 13524 18472 13530
rect 18420 13466 18472 13472
rect 18328 12912 18380 12918
rect 18234 12880 18290 12889
rect 18328 12854 18380 12860
rect 18234 12815 18290 12824
rect 18236 12776 18288 12782
rect 18236 12718 18288 12724
rect 18144 12368 18196 12374
rect 18144 12310 18196 12316
rect 17972 12260 18092 12288
rect 17696 12158 18000 12186
rect 17610 11996 17918 12005
rect 17610 11994 17616 11996
rect 17672 11994 17696 11996
rect 17752 11994 17776 11996
rect 17832 11994 17856 11996
rect 17912 11994 17918 11996
rect 17672 11942 17674 11994
rect 17854 11942 17856 11994
rect 17610 11940 17616 11942
rect 17672 11940 17696 11942
rect 17752 11940 17776 11942
rect 17832 11940 17856 11942
rect 17912 11940 17918 11942
rect 17610 11931 17918 11940
rect 17972 11778 18000 12158
rect 17880 11750 18000 11778
rect 17512 11614 17632 11642
rect 17500 11552 17552 11558
rect 17500 11494 17552 11500
rect 17512 11150 17540 11494
rect 17500 11144 17552 11150
rect 17500 11086 17552 11092
rect 17408 11076 17460 11082
rect 17408 11018 17460 11024
rect 17420 9654 17448 11018
rect 17604 10996 17632 11614
rect 17774 11248 17830 11257
rect 17774 11183 17830 11192
rect 17788 11150 17816 11183
rect 17776 11144 17828 11150
rect 17776 11086 17828 11092
rect 17880 11014 17908 11750
rect 17960 11280 18012 11286
rect 17958 11248 17960 11257
rect 18012 11248 18014 11257
rect 17958 11183 18014 11192
rect 18064 11150 18092 12260
rect 18144 12232 18196 12238
rect 18144 12174 18196 12180
rect 18156 12102 18184 12174
rect 18144 12096 18196 12102
rect 18144 12038 18196 12044
rect 18248 11830 18276 12718
rect 18512 12640 18564 12646
rect 18512 12582 18564 12588
rect 18524 12434 18552 12582
rect 18432 12406 18552 12434
rect 18236 11824 18288 11830
rect 18236 11766 18288 11772
rect 18326 11656 18382 11665
rect 18326 11591 18382 11600
rect 18052 11144 18104 11150
rect 18052 11086 18104 11092
rect 18142 11112 18198 11121
rect 18142 11047 18198 11056
rect 17512 10968 17632 10996
rect 17868 11008 17920 11014
rect 17512 10674 17540 10968
rect 17868 10950 17920 10956
rect 17610 10908 17918 10917
rect 17610 10906 17616 10908
rect 17672 10906 17696 10908
rect 17752 10906 17776 10908
rect 17832 10906 17856 10908
rect 17912 10906 17918 10908
rect 17672 10854 17674 10906
rect 17854 10854 17856 10906
rect 17610 10852 17616 10854
rect 17672 10852 17696 10854
rect 17752 10852 17776 10854
rect 17832 10852 17856 10854
rect 17912 10852 17918 10854
rect 17610 10843 17918 10852
rect 17776 10804 17828 10810
rect 17776 10746 17828 10752
rect 17788 10690 17816 10746
rect 17960 10736 18012 10742
rect 17500 10668 17552 10674
rect 17500 10610 17552 10616
rect 17696 10662 17816 10690
rect 17958 10704 17960 10713
rect 18012 10704 18014 10713
rect 17498 10568 17554 10577
rect 17498 10503 17500 10512
rect 17552 10503 17554 10512
rect 17500 10474 17552 10480
rect 17696 10130 17724 10662
rect 17958 10639 18014 10648
rect 18052 10668 18104 10674
rect 18052 10610 18104 10616
rect 17868 10464 17920 10470
rect 17868 10406 17920 10412
rect 17774 10160 17830 10169
rect 17684 10124 17736 10130
rect 17774 10095 17830 10104
rect 17684 10066 17736 10072
rect 17500 10056 17552 10062
rect 17498 10024 17500 10033
rect 17552 10024 17554 10033
rect 17788 9994 17816 10095
rect 17880 10010 17908 10406
rect 17498 9959 17554 9968
rect 17776 9988 17828 9994
rect 17880 9982 18000 10010
rect 17776 9930 17828 9936
rect 17500 9920 17552 9926
rect 17500 9862 17552 9868
rect 17408 9648 17460 9654
rect 17408 9590 17460 9596
rect 17512 9500 17540 9862
rect 17610 9820 17918 9829
rect 17610 9818 17616 9820
rect 17672 9818 17696 9820
rect 17752 9818 17776 9820
rect 17832 9818 17856 9820
rect 17912 9818 17918 9820
rect 17672 9766 17674 9818
rect 17854 9766 17856 9818
rect 17610 9764 17616 9766
rect 17672 9764 17696 9766
rect 17752 9764 17776 9766
rect 17832 9764 17856 9766
rect 17912 9764 17918 9766
rect 17610 9755 17918 9764
rect 17972 9704 18000 9982
rect 17420 9472 17540 9500
rect 17604 9676 18000 9704
rect 17316 5772 17368 5778
rect 17316 5714 17368 5720
rect 16764 5704 16816 5710
rect 16764 5646 16816 5652
rect 16776 5250 16804 5646
rect 16776 5222 16896 5250
rect 16672 5160 16724 5166
rect 16672 5102 16724 5108
rect 16764 5160 16816 5166
rect 16764 5102 16816 5108
rect 16672 5024 16724 5030
rect 16672 4966 16724 4972
rect 16580 3732 16632 3738
rect 16580 3674 16632 3680
rect 16580 3528 16632 3534
rect 16580 3470 16632 3476
rect 16592 3369 16620 3470
rect 16578 3360 16634 3369
rect 16578 3295 16634 3304
rect 16488 3052 16540 3058
rect 16488 2994 16540 3000
rect 16580 2440 16632 2446
rect 16580 2382 16632 2388
rect 16028 1080 16080 1086
rect 16028 1022 16080 1028
rect 15842 912 15898 921
rect 15476 876 15528 882
rect 15842 847 15898 856
rect 15476 818 15528 824
rect 16592 800 16620 2382
rect 16684 1737 16712 4966
rect 16670 1728 16726 1737
rect 16670 1663 16726 1672
rect 16776 1222 16804 5102
rect 16868 3534 16896 5222
rect 16950 4924 17258 4933
rect 16950 4922 16956 4924
rect 17012 4922 17036 4924
rect 17092 4922 17116 4924
rect 17172 4922 17196 4924
rect 17252 4922 17258 4924
rect 17012 4870 17014 4922
rect 17194 4870 17196 4922
rect 16950 4868 16956 4870
rect 17012 4868 17036 4870
rect 17092 4868 17116 4870
rect 17172 4868 17196 4870
rect 17252 4868 17258 4870
rect 16950 4859 17258 4868
rect 17316 4140 17368 4146
rect 17316 4082 17368 4088
rect 16950 3836 17258 3845
rect 16950 3834 16956 3836
rect 17012 3834 17036 3836
rect 17092 3834 17116 3836
rect 17172 3834 17196 3836
rect 17252 3834 17258 3836
rect 17012 3782 17014 3834
rect 17194 3782 17196 3834
rect 16950 3780 16956 3782
rect 17012 3780 17036 3782
rect 17092 3780 17116 3782
rect 17172 3780 17196 3782
rect 17252 3780 17258 3782
rect 16950 3771 17258 3780
rect 17328 3534 17356 4082
rect 17420 3942 17448 9472
rect 17604 8922 17632 9676
rect 17776 9580 17828 9586
rect 17776 9522 17828 9528
rect 17788 9382 17816 9522
rect 17776 9376 17828 9382
rect 17776 9318 17828 9324
rect 18064 8945 18092 10610
rect 18156 10470 18184 11047
rect 18144 10464 18196 10470
rect 18144 10406 18196 10412
rect 18156 10282 18184 10406
rect 18156 10254 18276 10282
rect 18142 10160 18198 10169
rect 18142 10095 18144 10104
rect 18196 10095 18198 10104
rect 18144 10066 18196 10072
rect 18144 9580 18196 9586
rect 18144 9522 18196 9528
rect 18156 9081 18184 9522
rect 18248 9178 18276 10254
rect 18236 9172 18288 9178
rect 18236 9114 18288 9120
rect 18142 9072 18198 9081
rect 18142 9007 18198 9016
rect 17512 8894 17632 8922
rect 18050 8936 18106 8945
rect 17512 6905 17540 8894
rect 18050 8871 18106 8880
rect 17960 8832 18012 8838
rect 17960 8774 18012 8780
rect 17610 8732 17918 8741
rect 17610 8730 17616 8732
rect 17672 8730 17696 8732
rect 17752 8730 17776 8732
rect 17832 8730 17856 8732
rect 17912 8730 17918 8732
rect 17672 8678 17674 8730
rect 17854 8678 17856 8730
rect 17610 8676 17616 8678
rect 17672 8676 17696 8678
rect 17752 8676 17776 8678
rect 17832 8676 17856 8678
rect 17912 8676 17918 8678
rect 17610 8667 17918 8676
rect 17592 8288 17644 8294
rect 17592 8230 17644 8236
rect 17604 7857 17632 8230
rect 17590 7848 17646 7857
rect 17590 7783 17646 7792
rect 17610 7644 17918 7653
rect 17610 7642 17616 7644
rect 17672 7642 17696 7644
rect 17752 7642 17776 7644
rect 17832 7642 17856 7644
rect 17912 7642 17918 7644
rect 17672 7590 17674 7642
rect 17854 7590 17856 7642
rect 17610 7588 17616 7590
rect 17672 7588 17696 7590
rect 17752 7588 17776 7590
rect 17832 7588 17856 7590
rect 17912 7588 17918 7590
rect 17610 7579 17918 7588
rect 17972 7274 18000 8774
rect 18052 8492 18104 8498
rect 18052 8434 18104 8440
rect 17960 7268 18012 7274
rect 17960 7210 18012 7216
rect 17498 6896 17554 6905
rect 17498 6831 17554 6840
rect 17500 6792 17552 6798
rect 17500 6734 17552 6740
rect 17512 5370 17540 6734
rect 17610 6556 17918 6565
rect 17610 6554 17616 6556
rect 17672 6554 17696 6556
rect 17752 6554 17776 6556
rect 17832 6554 17856 6556
rect 17912 6554 17918 6556
rect 17672 6502 17674 6554
rect 17854 6502 17856 6554
rect 17610 6500 17616 6502
rect 17672 6500 17696 6502
rect 17752 6500 17776 6502
rect 17832 6500 17856 6502
rect 17912 6500 17918 6502
rect 17610 6491 17918 6500
rect 17592 6452 17644 6458
rect 17592 6394 17644 6400
rect 17604 5710 17632 6394
rect 17960 6316 18012 6322
rect 17960 6258 18012 6264
rect 17972 5914 18000 6258
rect 17960 5908 18012 5914
rect 17960 5850 18012 5856
rect 17592 5704 17644 5710
rect 17592 5646 17644 5652
rect 17610 5468 17918 5477
rect 17610 5466 17616 5468
rect 17672 5466 17696 5468
rect 17752 5466 17776 5468
rect 17832 5466 17856 5468
rect 17912 5466 17918 5468
rect 17672 5414 17674 5466
rect 17854 5414 17856 5466
rect 17610 5412 17616 5414
rect 17672 5412 17696 5414
rect 17752 5412 17776 5414
rect 17832 5412 17856 5414
rect 17912 5412 17918 5414
rect 17610 5403 17918 5412
rect 17500 5364 17552 5370
rect 17500 5306 17552 5312
rect 17960 5228 18012 5234
rect 17960 5170 18012 5176
rect 17610 4380 17918 4389
rect 17610 4378 17616 4380
rect 17672 4378 17696 4380
rect 17752 4378 17776 4380
rect 17832 4378 17856 4380
rect 17912 4378 17918 4380
rect 17672 4326 17674 4378
rect 17854 4326 17856 4378
rect 17610 4324 17616 4326
rect 17672 4324 17696 4326
rect 17752 4324 17776 4326
rect 17832 4324 17856 4326
rect 17912 4324 17918 4326
rect 17610 4315 17918 4324
rect 17972 4078 18000 5170
rect 17960 4072 18012 4078
rect 17960 4014 18012 4020
rect 17868 4004 17920 4010
rect 17868 3946 17920 3952
rect 17408 3936 17460 3942
rect 17408 3878 17460 3884
rect 17880 3738 17908 3946
rect 17972 3738 18000 4014
rect 17868 3732 17920 3738
rect 17868 3674 17920 3680
rect 17960 3732 18012 3738
rect 17960 3674 18012 3680
rect 17958 3632 18014 3641
rect 17408 3596 17460 3602
rect 18064 3602 18092 8434
rect 18156 7886 18184 9007
rect 18144 7880 18196 7886
rect 18144 7822 18196 7828
rect 18340 5642 18368 11591
rect 18432 10810 18460 12406
rect 18604 12164 18656 12170
rect 18604 12106 18656 12112
rect 18512 11688 18564 11694
rect 18512 11630 18564 11636
rect 18420 10804 18472 10810
rect 18420 10746 18472 10752
rect 18420 10260 18472 10266
rect 18420 10202 18472 10208
rect 18432 9761 18460 10202
rect 18418 9752 18474 9761
rect 18418 9687 18474 9696
rect 18420 8832 18472 8838
rect 18418 8800 18420 8809
rect 18472 8800 18474 8809
rect 18418 8735 18474 8744
rect 18420 6656 18472 6662
rect 18420 6598 18472 6604
rect 18432 6361 18460 6598
rect 18418 6352 18474 6361
rect 18418 6287 18474 6296
rect 18328 5636 18380 5642
rect 18328 5578 18380 5584
rect 18326 5536 18382 5545
rect 18326 5471 18382 5480
rect 18340 5234 18368 5471
rect 18328 5228 18380 5234
rect 18328 5170 18380 5176
rect 18328 5024 18380 5030
rect 18328 4966 18380 4972
rect 18236 4140 18288 4146
rect 18236 4082 18288 4088
rect 18248 4049 18276 4082
rect 18234 4040 18290 4049
rect 18234 3975 18290 3984
rect 17958 3567 18014 3576
rect 18052 3596 18104 3602
rect 17408 3538 17460 3544
rect 16856 3528 16908 3534
rect 17316 3528 17368 3534
rect 16908 3488 16988 3516
rect 16856 3470 16908 3476
rect 16854 3360 16910 3369
rect 16854 3295 16910 3304
rect 16868 2854 16896 3295
rect 16960 2990 16988 3488
rect 17316 3470 17368 3476
rect 17420 3194 17448 3538
rect 17972 3534 18000 3567
rect 18052 3538 18104 3544
rect 17500 3528 17552 3534
rect 17500 3470 17552 3476
rect 17960 3528 18012 3534
rect 17960 3470 18012 3476
rect 17408 3188 17460 3194
rect 17408 3130 17460 3136
rect 16948 2984 17000 2990
rect 16948 2926 17000 2932
rect 17316 2984 17368 2990
rect 17316 2926 17368 2932
rect 16856 2848 16908 2854
rect 16856 2790 16908 2796
rect 16950 2748 17258 2757
rect 16950 2746 16956 2748
rect 17012 2746 17036 2748
rect 17092 2746 17116 2748
rect 17172 2746 17196 2748
rect 17252 2746 17258 2748
rect 17012 2694 17014 2746
rect 17194 2694 17196 2746
rect 16950 2692 16956 2694
rect 17012 2692 17036 2694
rect 17092 2692 17116 2694
rect 17172 2692 17196 2694
rect 17252 2692 17258 2694
rect 16950 2683 17258 2692
rect 16946 2544 17002 2553
rect 16946 2479 17002 2488
rect 16960 2446 16988 2479
rect 16948 2440 17000 2446
rect 16948 2382 17000 2388
rect 16856 2304 16908 2310
rect 16856 2246 16908 2252
rect 16868 2038 16896 2246
rect 16856 2032 16908 2038
rect 16856 1974 16908 1980
rect 16764 1216 16816 1222
rect 16764 1158 16816 1164
rect 17328 814 17356 2926
rect 17512 1562 17540 3470
rect 17610 3292 17918 3301
rect 17610 3290 17616 3292
rect 17672 3290 17696 3292
rect 17752 3290 17776 3292
rect 17832 3290 17856 3292
rect 17912 3290 17918 3292
rect 17672 3238 17674 3290
rect 17854 3238 17856 3290
rect 17610 3236 17616 3238
rect 17672 3236 17696 3238
rect 17752 3236 17776 3238
rect 17832 3236 17856 3238
rect 17912 3236 17918 3238
rect 17610 3227 17918 3236
rect 18064 2922 18092 3538
rect 18144 3528 18196 3534
rect 18142 3496 18144 3505
rect 18196 3496 18198 3505
rect 18142 3431 18198 3440
rect 18052 2916 18104 2922
rect 18052 2858 18104 2864
rect 18340 2530 18368 4966
rect 18420 3936 18472 3942
rect 18418 3904 18420 3913
rect 18472 3904 18474 3913
rect 18418 3839 18474 3848
rect 18248 2502 18368 2530
rect 18524 2514 18552 11630
rect 18616 8537 18644 12106
rect 18696 11008 18748 11014
rect 18696 10950 18748 10956
rect 18708 9110 18736 10950
rect 18696 9104 18748 9110
rect 18696 9046 18748 9052
rect 18800 8566 18828 15846
rect 18880 14272 18932 14278
rect 18880 14214 18932 14220
rect 18892 9994 18920 14214
rect 19340 13932 19392 13938
rect 19340 13874 19392 13880
rect 18972 12232 19024 12238
rect 18972 12174 19024 12180
rect 18880 9988 18932 9994
rect 18880 9930 18932 9936
rect 18788 8560 18840 8566
rect 18602 8528 18658 8537
rect 18788 8502 18840 8508
rect 18602 8463 18658 8472
rect 18892 8401 18920 9930
rect 18878 8392 18934 8401
rect 18878 8327 18934 8336
rect 18984 4486 19012 12174
rect 19248 12096 19300 12102
rect 19248 12038 19300 12044
rect 19156 10668 19208 10674
rect 19156 10610 19208 10616
rect 19064 10192 19116 10198
rect 19064 10134 19116 10140
rect 19076 7818 19104 10134
rect 19168 9489 19196 10610
rect 19154 9480 19210 9489
rect 19154 9415 19210 9424
rect 19064 7812 19116 7818
rect 19064 7754 19116 7760
rect 19260 6866 19288 12038
rect 19352 9586 19380 13874
rect 19432 13456 19484 13462
rect 19432 13398 19484 13404
rect 19340 9580 19392 9586
rect 19340 9522 19392 9528
rect 19248 6860 19300 6866
rect 19248 6802 19300 6808
rect 19444 6798 19472 13398
rect 19536 8430 19564 17750
rect 19524 8424 19576 8430
rect 19524 8366 19576 8372
rect 19432 6792 19484 6798
rect 19432 6734 19484 6740
rect 18972 4480 19024 4486
rect 18972 4422 19024 4428
rect 18512 2508 18564 2514
rect 17958 2408 18014 2417
rect 17958 2343 18014 2352
rect 17610 2204 17918 2213
rect 17610 2202 17616 2204
rect 17672 2202 17696 2204
rect 17752 2202 17776 2204
rect 17832 2202 17856 2204
rect 17912 2202 17918 2204
rect 17672 2150 17674 2202
rect 17854 2150 17856 2202
rect 17610 2148 17616 2150
rect 17672 2148 17696 2150
rect 17752 2148 17776 2150
rect 17832 2148 17856 2150
rect 17912 2148 17918 2150
rect 17610 2139 17918 2148
rect 17972 1902 18000 2343
rect 17960 1896 18012 1902
rect 17960 1838 18012 1844
rect 18248 1601 18276 2502
rect 18512 2450 18564 2456
rect 18328 2372 18380 2378
rect 18328 2314 18380 2320
rect 18234 1592 18290 1601
rect 17500 1556 17552 1562
rect 18234 1527 18290 1536
rect 17500 1498 17552 1504
rect 18340 1465 18368 2314
rect 18326 1456 18382 1465
rect 18326 1391 18382 1400
rect 17316 808 17368 814
rect 14648 536 14700 542
rect 14648 478 14700 484
rect 16578 0 16634 800
rect 17316 750 17368 756
<< via2 >>
rect 1122 18672 1178 18728
rect 754 17720 810 17776
rect 110 12280 166 12336
rect 386 6840 442 6896
rect 754 10104 810 10160
rect 754 9016 810 9072
rect 846 7248 902 7304
rect 1306 18264 1362 18320
rect 1490 16088 1546 16144
rect 2962 18536 3018 18592
rect 2318 17584 2374 17640
rect 1956 16890 2012 16892
rect 2036 16890 2092 16892
rect 2116 16890 2172 16892
rect 2196 16890 2252 16892
rect 1956 16838 2002 16890
rect 2002 16838 2012 16890
rect 2036 16838 2066 16890
rect 2066 16838 2078 16890
rect 2078 16838 2092 16890
rect 2116 16838 2130 16890
rect 2130 16838 2142 16890
rect 2142 16838 2172 16890
rect 2196 16838 2206 16890
rect 2206 16838 2252 16890
rect 1956 16836 2012 16838
rect 2036 16836 2092 16838
rect 2116 16836 2172 16838
rect 2196 16836 2252 16838
rect 1766 15952 1822 16008
rect 1582 15272 1638 15328
rect 1956 15802 2012 15804
rect 2036 15802 2092 15804
rect 2116 15802 2172 15804
rect 2196 15802 2252 15804
rect 1956 15750 2002 15802
rect 2002 15750 2012 15802
rect 2036 15750 2066 15802
rect 2066 15750 2078 15802
rect 2078 15750 2092 15802
rect 2116 15750 2130 15802
rect 2130 15750 2142 15802
rect 2142 15750 2172 15802
rect 2196 15750 2206 15802
rect 2206 15750 2252 15802
rect 1956 15748 2012 15750
rect 2036 15748 2092 15750
rect 2116 15748 2172 15750
rect 2196 15748 2252 15750
rect 1490 13640 1546 13696
rect 2616 17434 2672 17436
rect 2696 17434 2752 17436
rect 2776 17434 2832 17436
rect 2856 17434 2912 17436
rect 2616 17382 2662 17434
rect 2662 17382 2672 17434
rect 2696 17382 2726 17434
rect 2726 17382 2738 17434
rect 2738 17382 2752 17434
rect 2776 17382 2790 17434
rect 2790 17382 2802 17434
rect 2802 17382 2832 17434
rect 2856 17382 2866 17434
rect 2866 17382 2912 17434
rect 2616 17380 2672 17382
rect 2696 17380 2752 17382
rect 2776 17380 2832 17382
rect 2856 17380 2912 17382
rect 2410 16940 2412 16960
rect 2412 16940 2464 16960
rect 2464 16940 2466 16960
rect 2410 16904 2466 16940
rect 2616 16346 2672 16348
rect 2696 16346 2752 16348
rect 2776 16346 2832 16348
rect 2856 16346 2912 16348
rect 2616 16294 2662 16346
rect 2662 16294 2672 16346
rect 2696 16294 2726 16346
rect 2726 16294 2738 16346
rect 2738 16294 2752 16346
rect 2776 16294 2790 16346
rect 2790 16294 2802 16346
rect 2802 16294 2832 16346
rect 2856 16294 2866 16346
rect 2866 16294 2912 16346
rect 2616 16292 2672 16294
rect 2696 16292 2752 16294
rect 2776 16292 2832 16294
rect 2856 16292 2912 16294
rect 2502 15544 2558 15600
rect 1956 14714 2012 14716
rect 2036 14714 2092 14716
rect 2116 14714 2172 14716
rect 2196 14714 2252 14716
rect 1956 14662 2002 14714
rect 2002 14662 2012 14714
rect 2036 14662 2066 14714
rect 2066 14662 2078 14714
rect 2078 14662 2092 14714
rect 2116 14662 2130 14714
rect 2130 14662 2142 14714
rect 2142 14662 2172 14714
rect 2196 14662 2206 14714
rect 2206 14662 2252 14714
rect 1956 14660 2012 14662
rect 2036 14660 2092 14662
rect 2116 14660 2172 14662
rect 2196 14660 2252 14662
rect 1030 12392 1086 12448
rect 1214 12144 1270 12200
rect 1122 10920 1178 10976
rect 1030 9696 1086 9752
rect 1490 11600 1546 11656
rect 1398 11192 1454 11248
rect 1306 8336 1362 8392
rect 1858 14320 1914 14376
rect 2134 14184 2190 14240
rect 1950 13912 2006 13968
rect 1956 13626 2012 13628
rect 2036 13626 2092 13628
rect 2116 13626 2172 13628
rect 2196 13626 2252 13628
rect 1956 13574 2002 13626
rect 2002 13574 2012 13626
rect 2036 13574 2066 13626
rect 2066 13574 2078 13626
rect 2078 13574 2092 13626
rect 2116 13574 2130 13626
rect 2130 13574 2142 13626
rect 2142 13574 2172 13626
rect 2196 13574 2206 13626
rect 2206 13574 2252 13626
rect 1956 13572 2012 13574
rect 2036 13572 2092 13574
rect 2116 13572 2172 13574
rect 2196 13572 2252 13574
rect 1956 12538 2012 12540
rect 2036 12538 2092 12540
rect 2116 12538 2172 12540
rect 2196 12538 2252 12540
rect 1956 12486 2002 12538
rect 2002 12486 2012 12538
rect 2036 12486 2066 12538
rect 2066 12486 2078 12538
rect 2078 12486 2092 12538
rect 2116 12486 2130 12538
rect 2130 12486 2142 12538
rect 2142 12486 2172 12538
rect 2196 12486 2206 12538
rect 2206 12486 2252 12538
rect 1956 12484 2012 12486
rect 2036 12484 2092 12486
rect 2116 12484 2172 12486
rect 2196 12484 2252 12486
rect 2616 15258 2672 15260
rect 2696 15258 2752 15260
rect 2776 15258 2832 15260
rect 2856 15258 2912 15260
rect 2616 15206 2662 15258
rect 2662 15206 2672 15258
rect 2696 15206 2726 15258
rect 2726 15206 2738 15258
rect 2738 15206 2752 15258
rect 2776 15206 2790 15258
rect 2790 15206 2802 15258
rect 2802 15206 2832 15258
rect 2856 15206 2866 15258
rect 2866 15206 2912 15258
rect 2616 15204 2672 15206
rect 2696 15204 2752 15206
rect 2776 15204 2832 15206
rect 2856 15204 2912 15206
rect 2616 14170 2672 14172
rect 2696 14170 2752 14172
rect 2776 14170 2832 14172
rect 2856 14170 2912 14172
rect 2616 14118 2662 14170
rect 2662 14118 2672 14170
rect 2696 14118 2726 14170
rect 2726 14118 2738 14170
rect 2738 14118 2752 14170
rect 2776 14118 2790 14170
rect 2790 14118 2802 14170
rect 2802 14118 2832 14170
rect 2856 14118 2866 14170
rect 2866 14118 2912 14170
rect 2616 14116 2672 14118
rect 2696 14116 2752 14118
rect 2776 14116 2832 14118
rect 2856 14116 2912 14118
rect 2870 13268 2872 13288
rect 2872 13268 2924 13288
rect 2924 13268 2926 13288
rect 2870 13232 2926 13268
rect 2616 13082 2672 13084
rect 2696 13082 2752 13084
rect 2776 13082 2832 13084
rect 2856 13082 2912 13084
rect 2616 13030 2662 13082
rect 2662 13030 2672 13082
rect 2696 13030 2726 13082
rect 2726 13030 2738 13082
rect 2738 13030 2752 13082
rect 2776 13030 2790 13082
rect 2790 13030 2802 13082
rect 2802 13030 2832 13082
rect 2856 13030 2866 13082
rect 2866 13030 2912 13082
rect 2616 13028 2672 13030
rect 2696 13028 2752 13030
rect 2776 13028 2832 13030
rect 2856 13028 2912 13030
rect 1582 9016 1638 9072
rect 1490 6296 1546 6352
rect 1956 11450 2012 11452
rect 2036 11450 2092 11452
rect 2116 11450 2172 11452
rect 2196 11450 2252 11452
rect 1956 11398 2002 11450
rect 2002 11398 2012 11450
rect 2036 11398 2066 11450
rect 2066 11398 2078 11450
rect 2078 11398 2092 11450
rect 2116 11398 2130 11450
rect 2130 11398 2142 11450
rect 2142 11398 2172 11450
rect 2196 11398 2206 11450
rect 2206 11398 2252 11450
rect 1956 11396 2012 11398
rect 2036 11396 2092 11398
rect 2116 11396 2172 11398
rect 2196 11396 2252 11398
rect 1956 10362 2012 10364
rect 2036 10362 2092 10364
rect 2116 10362 2172 10364
rect 2196 10362 2252 10364
rect 1956 10310 2002 10362
rect 2002 10310 2012 10362
rect 2036 10310 2066 10362
rect 2066 10310 2078 10362
rect 2078 10310 2092 10362
rect 2116 10310 2130 10362
rect 2130 10310 2142 10362
rect 2142 10310 2172 10362
rect 2196 10310 2206 10362
rect 2206 10310 2252 10362
rect 1956 10308 2012 10310
rect 2036 10308 2092 10310
rect 2116 10308 2172 10310
rect 2196 10308 2252 10310
rect 2042 9424 2098 9480
rect 1956 9274 2012 9276
rect 2036 9274 2092 9276
rect 2116 9274 2172 9276
rect 2196 9274 2252 9276
rect 1956 9222 2002 9274
rect 2002 9222 2012 9274
rect 2036 9222 2066 9274
rect 2066 9222 2078 9274
rect 2078 9222 2092 9274
rect 2116 9222 2130 9274
rect 2130 9222 2142 9274
rect 2142 9222 2172 9274
rect 2196 9222 2206 9274
rect 2206 9222 2252 9274
rect 1956 9220 2012 9222
rect 2036 9220 2092 9222
rect 2116 9220 2172 9222
rect 2196 9220 2252 9222
rect 1214 3984 1270 4040
rect 938 3576 994 3632
rect 1398 4120 1454 4176
rect 1398 3848 1454 3904
rect 1766 7112 1822 7168
rect 1490 2352 1546 2408
rect 1950 8744 2006 8800
rect 2134 8880 2190 8936
rect 2226 8628 2282 8664
rect 2226 8608 2228 8628
rect 2228 8608 2280 8628
rect 2280 8608 2282 8628
rect 2594 12144 2650 12200
rect 2962 12824 3018 12880
rect 3146 14864 3202 14920
rect 2778 12688 2834 12744
rect 2870 12552 2926 12608
rect 2616 11994 2672 11996
rect 2696 11994 2752 11996
rect 2776 11994 2832 11996
rect 2856 11994 2912 11996
rect 2616 11942 2662 11994
rect 2662 11942 2672 11994
rect 2696 11942 2726 11994
rect 2726 11942 2738 11994
rect 2738 11942 2752 11994
rect 2776 11942 2790 11994
rect 2790 11942 2802 11994
rect 2802 11942 2832 11994
rect 2856 11942 2866 11994
rect 2866 11942 2912 11994
rect 2616 11940 2672 11942
rect 2696 11940 2752 11942
rect 2776 11940 2832 11942
rect 2856 11940 2912 11942
rect 2616 10906 2672 10908
rect 2696 10906 2752 10908
rect 2776 10906 2832 10908
rect 2856 10906 2912 10908
rect 2616 10854 2662 10906
rect 2662 10854 2672 10906
rect 2696 10854 2726 10906
rect 2726 10854 2738 10906
rect 2738 10854 2752 10906
rect 2776 10854 2790 10906
rect 2790 10854 2802 10906
rect 2802 10854 2832 10906
rect 2856 10854 2866 10906
rect 2866 10854 2912 10906
rect 2616 10852 2672 10854
rect 2696 10852 2752 10854
rect 2776 10852 2832 10854
rect 2856 10852 2912 10854
rect 2502 10648 2558 10704
rect 2410 9580 2466 9616
rect 2410 9560 2412 9580
rect 2412 9560 2464 9580
rect 2464 9560 2466 9580
rect 2778 10376 2834 10432
rect 2616 9818 2672 9820
rect 2696 9818 2752 9820
rect 2776 9818 2832 9820
rect 2856 9818 2912 9820
rect 2616 9766 2662 9818
rect 2662 9766 2672 9818
rect 2696 9766 2726 9818
rect 2726 9766 2738 9818
rect 2738 9766 2752 9818
rect 2776 9766 2790 9818
rect 2790 9766 2802 9818
rect 2802 9766 2832 9818
rect 2856 9766 2866 9818
rect 2866 9766 2912 9818
rect 2616 9764 2672 9766
rect 2696 9764 2752 9766
rect 2776 9764 2832 9766
rect 2856 9764 2912 9766
rect 2870 9596 2872 9616
rect 2872 9596 2924 9616
rect 2924 9596 2926 9616
rect 2870 9560 2926 9596
rect 3054 10512 3110 10568
rect 2594 9424 2650 9480
rect 2502 9016 2558 9072
rect 1956 8186 2012 8188
rect 2036 8186 2092 8188
rect 2116 8186 2172 8188
rect 2196 8186 2252 8188
rect 1956 8134 2002 8186
rect 2002 8134 2012 8186
rect 2036 8134 2066 8186
rect 2066 8134 2078 8186
rect 2078 8134 2092 8186
rect 2116 8134 2130 8186
rect 2130 8134 2142 8186
rect 2142 8134 2172 8186
rect 2196 8134 2206 8186
rect 2206 8134 2252 8186
rect 1956 8132 2012 8134
rect 2036 8132 2092 8134
rect 2116 8132 2172 8134
rect 2196 8132 2252 8134
rect 1956 7098 2012 7100
rect 2036 7098 2092 7100
rect 2116 7098 2172 7100
rect 2196 7098 2252 7100
rect 1956 7046 2002 7098
rect 2002 7046 2012 7098
rect 2036 7046 2066 7098
rect 2066 7046 2078 7098
rect 2078 7046 2092 7098
rect 2116 7046 2130 7098
rect 2130 7046 2142 7098
rect 2142 7046 2172 7098
rect 2196 7046 2206 7098
rect 2206 7046 2252 7098
rect 1956 7044 2012 7046
rect 2036 7044 2092 7046
rect 2116 7044 2172 7046
rect 2196 7044 2252 7046
rect 2226 6704 2282 6760
rect 2226 6160 2282 6216
rect 1956 6010 2012 6012
rect 2036 6010 2092 6012
rect 2116 6010 2172 6012
rect 2196 6010 2252 6012
rect 1956 5958 2002 6010
rect 2002 5958 2012 6010
rect 2036 5958 2066 6010
rect 2066 5958 2078 6010
rect 2078 5958 2092 6010
rect 2116 5958 2130 6010
rect 2130 5958 2142 6010
rect 2142 5958 2172 6010
rect 2196 5958 2206 6010
rect 2206 5958 2252 6010
rect 1956 5956 2012 5958
rect 2036 5956 2092 5958
rect 2116 5956 2172 5958
rect 2196 5956 2252 5958
rect 2962 9424 3018 9480
rect 3054 9288 3110 9344
rect 2962 9016 3018 9072
rect 2616 8730 2672 8732
rect 2696 8730 2752 8732
rect 2776 8730 2832 8732
rect 2856 8730 2912 8732
rect 2616 8678 2662 8730
rect 2662 8678 2672 8730
rect 2696 8678 2726 8730
rect 2726 8678 2738 8730
rect 2738 8678 2752 8730
rect 2776 8678 2790 8730
rect 2790 8678 2802 8730
rect 2802 8678 2832 8730
rect 2856 8678 2866 8730
rect 2866 8678 2912 8730
rect 2616 8676 2672 8678
rect 2696 8676 2752 8678
rect 2776 8676 2832 8678
rect 2856 8676 2912 8678
rect 2594 8472 2650 8528
rect 2616 7642 2672 7644
rect 2696 7642 2752 7644
rect 2776 7642 2832 7644
rect 2856 7642 2912 7644
rect 2616 7590 2662 7642
rect 2662 7590 2672 7642
rect 2696 7590 2726 7642
rect 2726 7590 2738 7642
rect 2738 7590 2752 7642
rect 2776 7590 2790 7642
rect 2790 7590 2802 7642
rect 2802 7590 2832 7642
rect 2856 7590 2866 7642
rect 2866 7590 2912 7642
rect 2616 7588 2672 7590
rect 2696 7588 2752 7590
rect 2776 7588 2832 7590
rect 2856 7588 2912 7590
rect 2410 6704 2466 6760
rect 2616 6554 2672 6556
rect 2696 6554 2752 6556
rect 2776 6554 2832 6556
rect 2856 6554 2912 6556
rect 2616 6502 2662 6554
rect 2662 6502 2672 6554
rect 2696 6502 2726 6554
rect 2726 6502 2738 6554
rect 2738 6502 2752 6554
rect 2776 6502 2790 6554
rect 2790 6502 2802 6554
rect 2802 6502 2832 6554
rect 2856 6502 2866 6554
rect 2866 6502 2912 6554
rect 2616 6500 2672 6502
rect 2696 6500 2752 6502
rect 2776 6500 2832 6502
rect 2856 6500 2912 6502
rect 1956 4922 2012 4924
rect 2036 4922 2092 4924
rect 2116 4922 2172 4924
rect 2196 4922 2252 4924
rect 1956 4870 2002 4922
rect 2002 4870 2012 4922
rect 2036 4870 2066 4922
rect 2066 4870 2078 4922
rect 2078 4870 2092 4922
rect 2116 4870 2130 4922
rect 2130 4870 2142 4922
rect 2142 4870 2172 4922
rect 2196 4870 2206 4922
rect 2206 4870 2252 4922
rect 1956 4868 2012 4870
rect 2036 4868 2092 4870
rect 2116 4868 2172 4870
rect 2196 4868 2252 4870
rect 2616 5466 2672 5468
rect 2696 5466 2752 5468
rect 2776 5466 2832 5468
rect 2856 5466 2912 5468
rect 2616 5414 2662 5466
rect 2662 5414 2672 5466
rect 2696 5414 2726 5466
rect 2726 5414 2738 5466
rect 2738 5414 2752 5466
rect 2776 5414 2790 5466
rect 2790 5414 2802 5466
rect 2802 5414 2832 5466
rect 2856 5414 2866 5466
rect 2866 5414 2912 5466
rect 2616 5412 2672 5414
rect 2696 5412 2752 5414
rect 2776 5412 2832 5414
rect 2856 5412 2912 5414
rect 2778 4800 2834 4856
rect 1956 3834 2012 3836
rect 2036 3834 2092 3836
rect 2116 3834 2172 3836
rect 2196 3834 2252 3836
rect 1956 3782 2002 3834
rect 2002 3782 2012 3834
rect 2036 3782 2066 3834
rect 2066 3782 2078 3834
rect 2078 3782 2092 3834
rect 2116 3782 2130 3834
rect 2130 3782 2142 3834
rect 2142 3782 2172 3834
rect 2196 3782 2206 3834
rect 2206 3782 2252 3834
rect 1956 3780 2012 3782
rect 2036 3780 2092 3782
rect 2116 3780 2172 3782
rect 2196 3780 2252 3782
rect 2616 4378 2672 4380
rect 2696 4378 2752 4380
rect 2776 4378 2832 4380
rect 2856 4378 2912 4380
rect 2616 4326 2662 4378
rect 2662 4326 2672 4378
rect 2696 4326 2726 4378
rect 2726 4326 2738 4378
rect 2738 4326 2752 4378
rect 2776 4326 2790 4378
rect 2790 4326 2802 4378
rect 2802 4326 2832 4378
rect 2856 4326 2866 4378
rect 2866 4326 2912 4378
rect 2616 4324 2672 4326
rect 2696 4324 2752 4326
rect 2776 4324 2832 4326
rect 2856 4324 2912 4326
rect 2410 3848 2466 3904
rect 1956 2746 2012 2748
rect 2036 2746 2092 2748
rect 2116 2746 2172 2748
rect 2196 2746 2252 2748
rect 1956 2694 2002 2746
rect 2002 2694 2012 2746
rect 2036 2694 2066 2746
rect 2066 2694 2078 2746
rect 2078 2694 2092 2746
rect 2116 2694 2130 2746
rect 2130 2694 2142 2746
rect 2142 2694 2172 2746
rect 2196 2694 2206 2746
rect 2206 2694 2252 2746
rect 1956 2692 2012 2694
rect 2036 2692 2092 2694
rect 2116 2692 2172 2694
rect 2196 2692 2252 2694
rect 3054 8064 3110 8120
rect 3238 12960 3294 13016
rect 3330 12824 3386 12880
rect 3054 5228 3110 5264
rect 3054 5208 3056 5228
rect 3056 5208 3108 5228
rect 3108 5208 3110 5228
rect 3054 3476 3056 3496
rect 3056 3476 3108 3496
rect 3108 3476 3110 3496
rect 3054 3440 3110 3476
rect 2616 3290 2672 3292
rect 2696 3290 2752 3292
rect 2776 3290 2832 3292
rect 2856 3290 2912 3292
rect 2616 3238 2662 3290
rect 2662 3238 2672 3290
rect 2696 3238 2726 3290
rect 2726 3238 2738 3290
rect 2738 3238 2752 3290
rect 2776 3238 2790 3290
rect 2790 3238 2802 3290
rect 2802 3238 2832 3290
rect 2856 3238 2866 3290
rect 2866 3238 2912 3290
rect 2616 3236 2672 3238
rect 2696 3236 2752 3238
rect 2776 3236 2832 3238
rect 2856 3236 2912 3238
rect 2778 3052 2834 3088
rect 4250 17856 4306 17912
rect 3882 17312 3938 17368
rect 3698 16224 3754 16280
rect 3422 12416 3478 12472
rect 4066 15564 4122 15600
rect 4066 15544 4068 15564
rect 4068 15544 4120 15564
rect 4120 15544 4122 15564
rect 4066 15408 4122 15464
rect 3882 12416 3938 12472
rect 3606 11872 3662 11928
rect 3514 10920 3570 10976
rect 3330 9696 3386 9752
rect 3330 9288 3386 9344
rect 3790 12008 3846 12064
rect 3514 10104 3570 10160
rect 3606 10004 3608 10024
rect 3608 10004 3660 10024
rect 3660 10004 3662 10024
rect 3606 9968 3662 10004
rect 3514 9868 3516 9888
rect 3516 9868 3568 9888
rect 3568 9868 3570 9888
rect 3514 9832 3570 9868
rect 3422 8744 3478 8800
rect 3606 9424 3662 9480
rect 3606 8744 3662 8800
rect 3514 8492 3570 8528
rect 3514 8472 3516 8492
rect 3516 8472 3568 8492
rect 3568 8472 3570 8492
rect 3514 8336 3570 8392
rect 3330 6432 3386 6488
rect 3606 8064 3662 8120
rect 4066 13504 4122 13560
rect 4250 13096 4306 13152
rect 4710 16088 4766 16144
rect 4434 14592 4490 14648
rect 4434 14456 4490 14512
rect 4342 12552 4398 12608
rect 4066 11736 4122 11792
rect 4250 11736 4306 11792
rect 3974 10376 4030 10432
rect 3974 10104 4030 10160
rect 3882 9288 3938 9344
rect 3882 8472 3938 8528
rect 4066 9288 4122 9344
rect 4526 14320 4582 14376
rect 4434 11328 4490 11384
rect 4894 15136 4950 15192
rect 4894 14220 4896 14240
rect 4896 14220 4948 14240
rect 4948 14220 4950 14240
rect 4894 14184 4950 14220
rect 4710 13776 4766 13832
rect 4618 12416 4674 12472
rect 4618 12280 4674 12336
rect 4802 11736 4858 11792
rect 4710 11328 4766 11384
rect 4618 11212 4674 11248
rect 4618 11192 4620 11212
rect 4620 11192 4672 11212
rect 4672 11192 4674 11212
rect 4342 9968 4398 10024
rect 4342 9696 4398 9752
rect 4158 8916 4160 8936
rect 4160 8916 4212 8936
rect 4212 8916 4214 8936
rect 3974 8064 4030 8120
rect 3790 7792 3846 7848
rect 3974 7384 4030 7440
rect 3882 6976 3938 7032
rect 3514 6160 3570 6216
rect 3514 5480 3570 5536
rect 3330 4256 3386 4312
rect 2778 3032 2780 3052
rect 2780 3032 2832 3052
rect 2832 3032 2834 3052
rect 3422 3304 3478 3360
rect 2410 1400 2466 1456
rect 2616 2202 2672 2204
rect 2696 2202 2752 2204
rect 2776 2202 2832 2204
rect 2856 2202 2912 2204
rect 2616 2150 2662 2202
rect 2662 2150 2672 2202
rect 2696 2150 2726 2202
rect 2726 2150 2738 2202
rect 2738 2150 2752 2202
rect 2776 2150 2790 2202
rect 2790 2150 2802 2202
rect 2802 2150 2832 2202
rect 2856 2150 2866 2202
rect 2866 2150 2912 2202
rect 2616 2148 2672 2150
rect 2696 2148 2752 2150
rect 2776 2148 2832 2150
rect 2856 2148 2912 2150
rect 2594 1400 2650 1456
rect 1398 992 1454 1048
rect 4158 8880 4214 8916
rect 4066 6840 4122 6896
rect 4158 6296 4214 6352
rect 3974 6180 4030 6216
rect 3974 6160 3976 6180
rect 3976 6160 4028 6180
rect 4028 6160 4030 6180
rect 3882 5752 3938 5808
rect 4066 5888 4122 5944
rect 3974 5344 4030 5400
rect 4986 13368 5042 13424
rect 5354 17176 5410 17232
rect 5446 16768 5502 16824
rect 5446 15000 5502 15056
rect 5814 17992 5870 18048
rect 5354 14048 5410 14104
rect 5446 13912 5502 13968
rect 5538 13504 5594 13560
rect 5630 12960 5686 13016
rect 5078 11328 5134 11384
rect 5078 11092 5080 11112
rect 5080 11092 5132 11112
rect 5132 11092 5134 11112
rect 5078 11056 5134 11092
rect 5354 11736 5410 11792
rect 5906 13776 5962 13832
rect 5814 13232 5870 13288
rect 5814 12280 5870 12336
rect 6366 18128 6422 18184
rect 6090 13504 6146 13560
rect 6550 16496 6606 16552
rect 6642 15272 6698 15328
rect 7616 17434 7672 17436
rect 7696 17434 7752 17436
rect 7776 17434 7832 17436
rect 7856 17434 7912 17436
rect 7616 17382 7662 17434
rect 7662 17382 7672 17434
rect 7696 17382 7726 17434
rect 7726 17382 7738 17434
rect 7738 17382 7752 17434
rect 7776 17382 7790 17434
rect 7790 17382 7802 17434
rect 7802 17382 7832 17434
rect 7856 17382 7866 17434
rect 7866 17382 7912 17434
rect 7616 17380 7672 17382
rect 7696 17380 7752 17382
rect 7776 17380 7832 17382
rect 7856 17380 7912 17382
rect 7470 17312 7526 17368
rect 6956 16890 7012 16892
rect 7036 16890 7092 16892
rect 7116 16890 7172 16892
rect 7196 16890 7252 16892
rect 6956 16838 7002 16890
rect 7002 16838 7012 16890
rect 7036 16838 7066 16890
rect 7066 16838 7078 16890
rect 7078 16838 7092 16890
rect 7116 16838 7130 16890
rect 7130 16838 7142 16890
rect 7142 16838 7172 16890
rect 7196 16838 7206 16890
rect 7206 16838 7252 16890
rect 6956 16836 7012 16838
rect 7036 16836 7092 16838
rect 7116 16836 7172 16838
rect 7196 16836 7252 16838
rect 7470 16768 7526 16824
rect 7616 16346 7672 16348
rect 7696 16346 7752 16348
rect 7776 16346 7832 16348
rect 7856 16346 7912 16348
rect 7616 16294 7662 16346
rect 7662 16294 7672 16346
rect 7696 16294 7726 16346
rect 7726 16294 7738 16346
rect 7738 16294 7752 16346
rect 7776 16294 7790 16346
rect 7790 16294 7802 16346
rect 7802 16294 7832 16346
rect 7856 16294 7866 16346
rect 7866 16294 7912 16346
rect 7616 16292 7672 16294
rect 7696 16292 7752 16294
rect 7776 16292 7832 16294
rect 7856 16292 7912 16294
rect 7470 16224 7526 16280
rect 7010 15952 7066 16008
rect 7378 15852 7380 15872
rect 7380 15852 7432 15872
rect 7432 15852 7434 15872
rect 7378 15816 7434 15852
rect 6956 15802 7012 15804
rect 7036 15802 7092 15804
rect 7116 15802 7172 15804
rect 7196 15802 7252 15804
rect 6956 15750 7002 15802
rect 7002 15750 7012 15802
rect 7036 15750 7066 15802
rect 7066 15750 7078 15802
rect 7078 15750 7092 15802
rect 7116 15750 7130 15802
rect 7130 15750 7142 15802
rect 7142 15750 7172 15802
rect 7196 15750 7206 15802
rect 7206 15750 7252 15802
rect 6956 15748 7012 15750
rect 7036 15748 7092 15750
rect 7116 15748 7172 15750
rect 7196 15748 7252 15750
rect 7470 15680 7526 15736
rect 6918 15544 6974 15600
rect 6956 14714 7012 14716
rect 7036 14714 7092 14716
rect 7116 14714 7172 14716
rect 7196 14714 7252 14716
rect 6956 14662 7002 14714
rect 7002 14662 7012 14714
rect 7036 14662 7066 14714
rect 7066 14662 7078 14714
rect 7078 14662 7092 14714
rect 7116 14662 7130 14714
rect 7130 14662 7142 14714
rect 7142 14662 7172 14714
rect 7196 14662 7206 14714
rect 7206 14662 7252 14714
rect 6956 14660 7012 14662
rect 7036 14660 7092 14662
rect 7116 14660 7172 14662
rect 7196 14660 7252 14662
rect 6458 13776 6514 13832
rect 6458 13504 6514 13560
rect 6182 13232 6238 13288
rect 6182 12824 6238 12880
rect 5998 11736 6054 11792
rect 5722 11328 5778 11384
rect 5906 11600 5962 11656
rect 5814 11192 5870 11248
rect 4986 10104 5042 10160
rect 4802 9560 4858 9616
rect 4894 9424 4950 9480
rect 4618 8200 4674 8256
rect 4434 6568 4490 6624
rect 3974 4936 4030 4992
rect 3882 3984 3938 4040
rect 3238 2080 3294 2136
rect 4710 7248 4766 7304
rect 4894 8200 4950 8256
rect 4342 3848 4398 3904
rect 4894 6568 4950 6624
rect 4894 6160 4950 6216
rect 5446 10648 5502 10704
rect 5262 9696 5318 9752
rect 5170 9460 5172 9480
rect 5172 9460 5224 9480
rect 5224 9460 5226 9480
rect 5170 9424 5226 9460
rect 5078 8336 5134 8392
rect 4802 4664 4858 4720
rect 4710 4548 4766 4584
rect 4710 4528 4712 4548
rect 4712 4528 4764 4548
rect 4764 4528 4766 4548
rect 4618 3712 4674 3768
rect 4526 3476 4528 3496
rect 4528 3476 4580 3496
rect 4580 3476 4582 3496
rect 4526 3440 4582 3476
rect 5354 8916 5356 8936
rect 5356 8916 5408 8936
rect 5408 8916 5410 8936
rect 5354 8880 5410 8916
rect 5262 8744 5318 8800
rect 5262 8472 5318 8528
rect 5262 8084 5318 8120
rect 5262 8064 5264 8084
rect 5264 8064 5316 8084
rect 5316 8064 5318 8084
rect 5170 5072 5226 5128
rect 4986 3984 5042 4040
rect 4986 3848 5042 3904
rect 4986 3032 5042 3088
rect 4802 1128 4858 1184
rect 6182 11464 6238 11520
rect 6182 10920 6238 10976
rect 6366 12960 6422 13016
rect 7286 13912 7342 13968
rect 6366 12552 6422 12608
rect 6366 12144 6422 12200
rect 6550 12844 6606 12880
rect 6550 12824 6552 12844
rect 6552 12824 6604 12844
rect 6604 12824 6606 12844
rect 6550 12688 6606 12744
rect 5998 10532 6054 10568
rect 5998 10512 6000 10532
rect 6000 10512 6052 10532
rect 6052 10512 6054 10532
rect 6090 9968 6146 10024
rect 5722 6840 5778 6896
rect 5814 5888 5870 5944
rect 5722 5208 5778 5264
rect 5446 4528 5502 4584
rect 5446 4120 5502 4176
rect 5998 9152 6054 9208
rect 5998 8372 6000 8392
rect 6000 8372 6052 8392
rect 6052 8372 6054 8392
rect 5998 8336 6054 8372
rect 6274 10784 6330 10840
rect 6458 10920 6514 10976
rect 6458 10648 6514 10704
rect 6458 10512 6514 10568
rect 6090 6704 6146 6760
rect 6458 9968 6514 10024
rect 6458 9696 6514 9752
rect 6366 9288 6422 9344
rect 6274 6704 6330 6760
rect 5446 3576 5502 3632
rect 5630 3440 5686 3496
rect 5538 3304 5594 3360
rect 5814 4392 5870 4448
rect 5906 3884 5908 3904
rect 5908 3884 5960 3904
rect 5960 3884 5962 3904
rect 5906 3848 5962 3884
rect 6090 4256 6146 4312
rect 6090 3476 6092 3496
rect 6092 3476 6144 3496
rect 6144 3476 6146 3496
rect 6090 3440 6146 3476
rect 6090 1808 6146 1864
rect 6274 6160 6330 6216
rect 6458 7520 6514 7576
rect 6734 12688 6790 12744
rect 6956 13626 7012 13628
rect 7036 13626 7092 13628
rect 7116 13626 7172 13628
rect 7196 13626 7252 13628
rect 6956 13574 7002 13626
rect 7002 13574 7012 13626
rect 7036 13574 7066 13626
rect 7066 13574 7078 13626
rect 7078 13574 7092 13626
rect 7116 13574 7130 13626
rect 7130 13574 7142 13626
rect 7142 13574 7172 13626
rect 7196 13574 7206 13626
rect 7206 13574 7252 13626
rect 6956 13572 7012 13574
rect 7036 13572 7092 13574
rect 7116 13572 7172 13574
rect 7196 13572 7252 13574
rect 7194 13232 7250 13288
rect 7378 13096 7434 13152
rect 7286 12960 7342 13016
rect 7616 15258 7672 15260
rect 7696 15258 7752 15260
rect 7776 15258 7832 15260
rect 7856 15258 7912 15260
rect 7616 15206 7662 15258
rect 7662 15206 7672 15258
rect 7696 15206 7726 15258
rect 7726 15206 7738 15258
rect 7738 15206 7752 15258
rect 7776 15206 7790 15258
rect 7790 15206 7802 15258
rect 7802 15206 7832 15258
rect 7856 15206 7866 15258
rect 7866 15206 7912 15258
rect 7616 15204 7672 15206
rect 7696 15204 7752 15206
rect 7776 15204 7832 15206
rect 7856 15204 7912 15206
rect 7616 14170 7672 14172
rect 7696 14170 7752 14172
rect 7776 14170 7832 14172
rect 7856 14170 7912 14172
rect 7616 14118 7662 14170
rect 7662 14118 7672 14170
rect 7696 14118 7726 14170
rect 7726 14118 7738 14170
rect 7738 14118 7752 14170
rect 7776 14118 7790 14170
rect 7790 14118 7802 14170
rect 7802 14118 7832 14170
rect 7856 14118 7866 14170
rect 7866 14118 7912 14170
rect 7616 14116 7672 14118
rect 7696 14116 7752 14118
rect 7776 14116 7832 14118
rect 7856 14116 7912 14118
rect 8666 17040 8722 17096
rect 8206 14592 8262 14648
rect 8482 15136 8538 15192
rect 8298 14320 8354 14376
rect 7930 13504 7986 13560
rect 7562 13232 7618 13288
rect 7746 13232 7802 13288
rect 7616 13082 7672 13084
rect 7696 13082 7752 13084
rect 7776 13082 7832 13084
rect 7856 13082 7912 13084
rect 7616 13030 7662 13082
rect 7662 13030 7672 13082
rect 7696 13030 7726 13082
rect 7726 13030 7738 13082
rect 7738 13030 7752 13082
rect 7776 13030 7790 13082
rect 7790 13030 7802 13082
rect 7802 13030 7832 13082
rect 7856 13030 7866 13082
rect 7866 13030 7912 13082
rect 7616 13028 7672 13030
rect 7696 13028 7752 13030
rect 7776 13028 7832 13030
rect 7856 13028 7912 13030
rect 6956 12538 7012 12540
rect 7036 12538 7092 12540
rect 7116 12538 7172 12540
rect 7196 12538 7252 12540
rect 6956 12486 7002 12538
rect 7002 12486 7012 12538
rect 7036 12486 7066 12538
rect 7066 12486 7078 12538
rect 7078 12486 7092 12538
rect 7116 12486 7130 12538
rect 7130 12486 7142 12538
rect 7142 12486 7172 12538
rect 7196 12486 7206 12538
rect 7206 12486 7252 12538
rect 6956 12484 7012 12486
rect 7036 12484 7092 12486
rect 7116 12484 7172 12486
rect 7196 12484 7252 12486
rect 7470 12552 7526 12608
rect 7654 12280 7710 12336
rect 7102 12144 7158 12200
rect 6734 11464 6790 11520
rect 7102 11600 7158 11656
rect 8298 13368 8354 13424
rect 9126 17176 9182 17232
rect 9126 16632 9182 16688
rect 8942 15408 8998 15464
rect 9126 15408 9182 15464
rect 8850 15272 8906 15328
rect 8574 13912 8630 13968
rect 8574 13232 8630 13288
rect 8482 13096 8538 13152
rect 7616 11994 7672 11996
rect 7696 11994 7752 11996
rect 7776 11994 7832 11996
rect 7856 11994 7912 11996
rect 7616 11942 7662 11994
rect 7662 11942 7672 11994
rect 7696 11942 7726 11994
rect 7726 11942 7738 11994
rect 7738 11942 7752 11994
rect 7776 11942 7790 11994
rect 7790 11942 7802 11994
rect 7802 11942 7832 11994
rect 7856 11942 7866 11994
rect 7866 11942 7912 11994
rect 7616 11940 7672 11942
rect 7696 11940 7752 11942
rect 7776 11940 7832 11942
rect 7856 11940 7912 11942
rect 8022 11872 8078 11928
rect 7378 11464 7434 11520
rect 6956 11450 7012 11452
rect 7036 11450 7092 11452
rect 7116 11450 7172 11452
rect 7196 11450 7252 11452
rect 6956 11398 7002 11450
rect 7002 11398 7012 11450
rect 7036 11398 7066 11450
rect 7066 11398 7078 11450
rect 7078 11398 7092 11450
rect 7116 11398 7130 11450
rect 7130 11398 7142 11450
rect 7142 11398 7172 11450
rect 7196 11398 7206 11450
rect 7206 11398 7252 11450
rect 6956 11396 7012 11398
rect 7036 11396 7092 11398
rect 7116 11396 7172 11398
rect 7196 11396 7252 11398
rect 6918 10920 6974 10976
rect 6826 10784 6882 10840
rect 7010 10648 7066 10704
rect 7286 10920 7342 10976
rect 7930 11328 7986 11384
rect 7930 11192 7986 11248
rect 7616 10906 7672 10908
rect 7696 10906 7752 10908
rect 7776 10906 7832 10908
rect 7856 10906 7912 10908
rect 7616 10854 7662 10906
rect 7662 10854 7672 10906
rect 7696 10854 7726 10906
rect 7726 10854 7738 10906
rect 7738 10854 7752 10906
rect 7776 10854 7790 10906
rect 7790 10854 7802 10906
rect 7802 10854 7832 10906
rect 7856 10854 7866 10906
rect 7866 10854 7912 10906
rect 7616 10852 7672 10854
rect 7696 10852 7752 10854
rect 7776 10852 7832 10854
rect 7856 10852 7912 10854
rect 7470 10648 7526 10704
rect 6956 10362 7012 10364
rect 7036 10362 7092 10364
rect 7116 10362 7172 10364
rect 7196 10362 7252 10364
rect 6956 10310 7002 10362
rect 7002 10310 7012 10362
rect 7036 10310 7066 10362
rect 7066 10310 7078 10362
rect 7078 10310 7092 10362
rect 7116 10310 7130 10362
rect 7130 10310 7142 10362
rect 7142 10310 7172 10362
rect 7196 10310 7206 10362
rect 7206 10310 7252 10362
rect 6956 10308 7012 10310
rect 7036 10308 7092 10310
rect 7116 10308 7172 10310
rect 7196 10308 7252 10310
rect 7470 10376 7526 10432
rect 7654 10240 7710 10296
rect 6956 9274 7012 9276
rect 7036 9274 7092 9276
rect 7116 9274 7172 9276
rect 7196 9274 7252 9276
rect 6956 9222 7002 9274
rect 7002 9222 7012 9274
rect 7036 9222 7066 9274
rect 7066 9222 7078 9274
rect 7078 9222 7092 9274
rect 7116 9222 7130 9274
rect 7130 9222 7142 9274
rect 7142 9222 7172 9274
rect 7196 9222 7206 9274
rect 7206 9222 7252 9274
rect 6956 9220 7012 9222
rect 7036 9220 7092 9222
rect 7116 9220 7172 9222
rect 7196 9220 7252 9222
rect 7010 8608 7066 8664
rect 6642 8200 6698 8256
rect 6734 8064 6790 8120
rect 7378 9288 7434 9344
rect 7378 9152 7434 9208
rect 7378 8880 7434 8936
rect 7378 8744 7434 8800
rect 7286 8472 7342 8528
rect 6956 8186 7012 8188
rect 7036 8186 7092 8188
rect 7116 8186 7172 8188
rect 7196 8186 7252 8188
rect 6956 8134 7002 8186
rect 7002 8134 7012 8186
rect 7036 8134 7066 8186
rect 7066 8134 7078 8186
rect 7078 8134 7092 8186
rect 7116 8134 7130 8186
rect 7130 8134 7142 8186
rect 7142 8134 7172 8186
rect 7196 8134 7206 8186
rect 7206 8134 7252 8186
rect 6956 8132 7012 8134
rect 7036 8132 7092 8134
rect 7116 8132 7172 8134
rect 7196 8132 7252 8134
rect 6458 5752 6514 5808
rect 6458 3712 6514 3768
rect 6642 6740 6644 6760
rect 6644 6740 6696 6760
rect 6696 6740 6698 6760
rect 6642 6704 6698 6740
rect 6642 6160 6698 6216
rect 7102 7928 7158 7984
rect 7194 7656 7250 7712
rect 6956 7098 7012 7100
rect 7036 7098 7092 7100
rect 7116 7098 7172 7100
rect 7196 7098 7252 7100
rect 6956 7046 7002 7098
rect 7002 7046 7012 7098
rect 7036 7046 7066 7098
rect 7066 7046 7078 7098
rect 7078 7046 7092 7098
rect 7116 7046 7130 7098
rect 7130 7046 7142 7098
rect 7142 7046 7172 7098
rect 7196 7046 7206 7098
rect 7206 7046 7252 7098
rect 6956 7044 7012 7046
rect 7036 7044 7092 7046
rect 7116 7044 7172 7046
rect 7196 7044 7252 7046
rect 7378 6568 7434 6624
rect 7286 6432 7342 6488
rect 6956 6010 7012 6012
rect 7036 6010 7092 6012
rect 7116 6010 7172 6012
rect 7196 6010 7252 6012
rect 6956 5958 7002 6010
rect 7002 5958 7012 6010
rect 7036 5958 7066 6010
rect 7066 5958 7078 6010
rect 7078 5958 7092 6010
rect 7116 5958 7130 6010
rect 7130 5958 7142 6010
rect 7142 5958 7172 6010
rect 7196 5958 7206 6010
rect 7206 5958 7252 6010
rect 6956 5956 7012 5958
rect 7036 5956 7092 5958
rect 7116 5956 7172 5958
rect 7196 5956 7252 5958
rect 7010 5752 7066 5808
rect 6734 5516 6736 5536
rect 6736 5516 6788 5536
rect 6788 5516 6790 5536
rect 6734 5480 6790 5516
rect 6734 4972 6736 4992
rect 6736 4972 6788 4992
rect 6788 4972 6790 4992
rect 6734 4936 6790 4972
rect 6642 4664 6698 4720
rect 6642 4392 6698 4448
rect 7102 5616 7158 5672
rect 7286 5480 7342 5536
rect 6956 4922 7012 4924
rect 7036 4922 7092 4924
rect 7116 4922 7172 4924
rect 7196 4922 7252 4924
rect 6956 4870 7002 4922
rect 7002 4870 7012 4922
rect 7036 4870 7066 4922
rect 7066 4870 7078 4922
rect 7078 4870 7092 4922
rect 7116 4870 7130 4922
rect 7130 4870 7142 4922
rect 7142 4870 7172 4922
rect 7196 4870 7206 4922
rect 7206 4870 7252 4922
rect 6956 4868 7012 4870
rect 7036 4868 7092 4870
rect 7116 4868 7172 4870
rect 7196 4868 7252 4870
rect 7194 4120 7250 4176
rect 6956 3834 7012 3836
rect 7036 3834 7092 3836
rect 7116 3834 7172 3836
rect 7196 3834 7252 3836
rect 6956 3782 7002 3834
rect 7002 3782 7012 3834
rect 7036 3782 7066 3834
rect 7066 3782 7078 3834
rect 7078 3782 7092 3834
rect 7116 3782 7130 3834
rect 7130 3782 7142 3834
rect 7142 3782 7172 3834
rect 7196 3782 7206 3834
rect 7206 3782 7252 3834
rect 6956 3780 7012 3782
rect 7036 3780 7092 3782
rect 7116 3780 7172 3782
rect 7196 3780 7252 3782
rect 7010 3576 7066 3632
rect 7194 3576 7250 3632
rect 7616 9818 7672 9820
rect 7696 9818 7752 9820
rect 7776 9818 7832 9820
rect 7856 9818 7912 9820
rect 7616 9766 7662 9818
rect 7662 9766 7672 9818
rect 7696 9766 7726 9818
rect 7726 9766 7738 9818
rect 7738 9766 7752 9818
rect 7776 9766 7790 9818
rect 7790 9766 7802 9818
rect 7802 9766 7832 9818
rect 7856 9766 7866 9818
rect 7866 9766 7912 9818
rect 7616 9764 7672 9766
rect 7696 9764 7752 9766
rect 7776 9764 7832 9766
rect 7856 9764 7912 9766
rect 7654 8880 7710 8936
rect 8206 10260 8262 10296
rect 8206 10240 8208 10260
rect 8208 10240 8260 10260
rect 8260 10240 8262 10260
rect 8206 9832 8262 9888
rect 7616 8730 7672 8732
rect 7696 8730 7752 8732
rect 7776 8730 7832 8732
rect 7856 8730 7912 8732
rect 7616 8678 7662 8730
rect 7662 8678 7672 8730
rect 7696 8678 7726 8730
rect 7726 8678 7738 8730
rect 7738 8678 7752 8730
rect 7776 8678 7790 8730
rect 7790 8678 7802 8730
rect 7802 8678 7832 8730
rect 7856 8678 7866 8730
rect 7866 8678 7912 8730
rect 7616 8676 7672 8678
rect 7696 8676 7752 8678
rect 7776 8676 7832 8678
rect 7856 8676 7912 8678
rect 7562 8200 7618 8256
rect 7562 8064 7618 8120
rect 7746 7928 7802 7984
rect 7930 8200 7986 8256
rect 7616 7642 7672 7644
rect 7696 7642 7752 7644
rect 7776 7642 7832 7644
rect 7856 7642 7912 7644
rect 7616 7590 7662 7642
rect 7662 7590 7672 7642
rect 7696 7590 7726 7642
rect 7726 7590 7738 7642
rect 7738 7590 7752 7642
rect 7776 7590 7790 7642
rect 7790 7590 7802 7642
rect 7802 7590 7832 7642
rect 7856 7590 7866 7642
rect 7866 7590 7912 7642
rect 7616 7588 7672 7590
rect 7696 7588 7752 7590
rect 7776 7588 7832 7590
rect 7856 7588 7912 7590
rect 7562 7248 7618 7304
rect 8114 9036 8170 9072
rect 8114 9016 8116 9036
rect 8116 9016 8168 9036
rect 8168 9016 8170 9036
rect 8114 7928 8170 7984
rect 8298 8744 8354 8800
rect 8390 8608 8446 8664
rect 8298 7928 8354 7984
rect 7562 6740 7564 6760
rect 7564 6740 7616 6760
rect 7616 6740 7618 6760
rect 7562 6704 7618 6740
rect 8298 7112 8354 7168
rect 7616 6554 7672 6556
rect 7696 6554 7752 6556
rect 7776 6554 7832 6556
rect 7856 6554 7912 6556
rect 7616 6502 7662 6554
rect 7662 6502 7672 6554
rect 7696 6502 7726 6554
rect 7726 6502 7738 6554
rect 7738 6502 7752 6554
rect 7776 6502 7790 6554
rect 7790 6502 7802 6554
rect 7802 6502 7832 6554
rect 7856 6502 7866 6554
rect 7866 6502 7912 6554
rect 7616 6500 7672 6502
rect 7696 6500 7752 6502
rect 7776 6500 7832 6502
rect 7856 6500 7912 6502
rect 7654 5888 7710 5944
rect 8022 6024 8078 6080
rect 7616 5466 7672 5468
rect 7696 5466 7752 5468
rect 7776 5466 7832 5468
rect 7856 5466 7912 5468
rect 7616 5414 7662 5466
rect 7662 5414 7672 5466
rect 7696 5414 7726 5466
rect 7726 5414 7738 5466
rect 7738 5414 7752 5466
rect 7776 5414 7790 5466
rect 7790 5414 7802 5466
rect 7802 5414 7832 5466
rect 7856 5414 7866 5466
rect 7866 5414 7912 5466
rect 7616 5412 7672 5414
rect 7696 5412 7752 5414
rect 7776 5412 7832 5414
rect 7856 5412 7912 5414
rect 7470 5364 7526 5400
rect 7470 5344 7472 5364
rect 7472 5344 7524 5364
rect 7524 5344 7526 5364
rect 7378 4256 7434 4312
rect 7930 4528 7986 4584
rect 7616 4378 7672 4380
rect 7696 4378 7752 4380
rect 7776 4378 7832 4380
rect 7856 4378 7912 4380
rect 7616 4326 7662 4378
rect 7662 4326 7672 4378
rect 7696 4326 7726 4378
rect 7726 4326 7738 4378
rect 7738 4326 7752 4378
rect 7776 4326 7790 4378
rect 7790 4326 7802 4378
rect 7802 4326 7832 4378
rect 7856 4326 7866 4378
rect 7866 4326 7912 4378
rect 7616 4324 7672 4326
rect 7696 4324 7752 4326
rect 7776 4324 7832 4326
rect 7856 4324 7912 4326
rect 8390 5344 8446 5400
rect 8390 4392 8446 4448
rect 8390 3984 8446 4040
rect 8206 3576 8262 3632
rect 7286 3304 7342 3360
rect 6550 2624 6606 2680
rect 6550 1536 6606 1592
rect 6956 2746 7012 2748
rect 7036 2746 7092 2748
rect 7116 2746 7172 2748
rect 7196 2746 7252 2748
rect 6956 2694 7002 2746
rect 7002 2694 7012 2746
rect 7036 2694 7066 2746
rect 7066 2694 7078 2746
rect 7078 2694 7092 2746
rect 7116 2694 7130 2746
rect 7130 2694 7142 2746
rect 7142 2694 7172 2746
rect 7196 2694 7206 2746
rect 7206 2694 7252 2746
rect 6956 2692 7012 2694
rect 7036 2692 7092 2694
rect 7116 2692 7172 2694
rect 7196 2692 7252 2694
rect 7194 1400 7250 1456
rect 7616 3290 7672 3292
rect 7696 3290 7752 3292
rect 7776 3290 7832 3292
rect 7856 3290 7912 3292
rect 7616 3238 7662 3290
rect 7662 3238 7672 3290
rect 7696 3238 7726 3290
rect 7726 3238 7738 3290
rect 7738 3238 7752 3290
rect 7776 3238 7790 3290
rect 7790 3238 7802 3290
rect 7802 3238 7832 3290
rect 7856 3238 7866 3290
rect 7866 3238 7912 3290
rect 7616 3236 7672 3238
rect 7696 3236 7752 3238
rect 7776 3236 7832 3238
rect 7856 3236 7912 3238
rect 7930 2932 7932 2952
rect 7932 2932 7984 2952
rect 7984 2932 7986 2952
rect 7930 2896 7986 2932
rect 8298 3168 8354 3224
rect 8574 10512 8630 10568
rect 9310 14320 9366 14376
rect 9034 9288 9090 9344
rect 9218 13232 9274 13288
rect 9310 13096 9366 13152
rect 9218 11328 9274 11384
rect 9218 8880 9274 8936
rect 8574 3848 8630 3904
rect 8298 2896 8354 2952
rect 8206 2624 8262 2680
rect 7470 2216 7526 2272
rect 8022 2216 8078 2272
rect 7616 2202 7672 2204
rect 7696 2202 7752 2204
rect 7776 2202 7832 2204
rect 7856 2202 7912 2204
rect 7616 2150 7662 2202
rect 7662 2150 7672 2202
rect 7696 2150 7726 2202
rect 7726 2150 7738 2202
rect 7738 2150 7752 2202
rect 7776 2150 7790 2202
rect 7790 2150 7802 2202
rect 7802 2150 7832 2202
rect 7856 2150 7866 2202
rect 7866 2150 7912 2202
rect 7616 2148 7672 2150
rect 7696 2148 7752 2150
rect 7776 2148 7832 2150
rect 7856 2148 7912 2150
rect 9034 6704 9090 6760
rect 8942 6568 8998 6624
rect 8942 5908 8998 5944
rect 8942 5888 8944 5908
rect 8944 5888 8996 5908
rect 8996 5888 8998 5908
rect 8850 5244 8852 5264
rect 8852 5244 8904 5264
rect 8904 5244 8906 5264
rect 8850 5208 8906 5244
rect 9126 5516 9128 5536
rect 9128 5516 9180 5536
rect 9180 5516 9182 5536
rect 9126 5480 9182 5516
rect 8850 4392 8906 4448
rect 8850 3984 8906 4040
rect 8666 2624 8722 2680
rect 8574 2508 8630 2544
rect 8574 2488 8576 2508
rect 8576 2488 8628 2508
rect 8628 2488 8630 2508
rect 8942 3848 8998 3904
rect 9862 16496 9918 16552
rect 9770 15020 9826 15056
rect 9770 15000 9772 15020
rect 9772 15000 9824 15020
rect 9824 15000 9826 15020
rect 9770 14320 9826 14376
rect 9862 12960 9918 13016
rect 9678 12824 9734 12880
rect 10874 18536 10930 18592
rect 10138 13368 10194 13424
rect 9770 12724 9772 12744
rect 9772 12724 9824 12744
rect 9824 12724 9826 12744
rect 9770 12688 9826 12724
rect 10138 12824 10194 12880
rect 9954 12552 10010 12608
rect 9678 12008 9734 12064
rect 9494 10240 9550 10296
rect 9770 11600 9826 11656
rect 9678 11464 9734 11520
rect 9678 11192 9734 11248
rect 9494 9832 9550 9888
rect 9310 7112 9366 7168
rect 9770 10920 9826 10976
rect 9954 12144 10010 12200
rect 10598 16224 10654 16280
rect 12346 17856 12402 17912
rect 11518 16904 11574 16960
rect 11334 16632 11390 16688
rect 10598 15700 10654 15736
rect 10598 15680 10600 15700
rect 10600 15680 10652 15700
rect 10652 15680 10654 15700
rect 10598 15444 10600 15464
rect 10600 15444 10652 15464
rect 10652 15444 10654 15464
rect 10598 15408 10654 15444
rect 10506 15000 10562 15056
rect 10506 13912 10562 13968
rect 10414 13776 10470 13832
rect 9954 11464 10010 11520
rect 9954 10784 10010 10840
rect 9862 9424 9918 9480
rect 9770 8744 9826 8800
rect 9770 8472 9826 8528
rect 9586 8064 9642 8120
rect 9770 8200 9826 8256
rect 9494 7656 9550 7712
rect 9678 7656 9734 7712
rect 9586 6704 9642 6760
rect 9586 6432 9642 6488
rect 9494 5752 9550 5808
rect 9678 6316 9734 6352
rect 9678 6296 9680 6316
rect 9680 6296 9732 6316
rect 9732 6296 9734 6316
rect 10230 10240 10286 10296
rect 10598 12824 10654 12880
rect 10874 14728 10930 14784
rect 10966 14456 11022 14512
rect 11242 14592 11298 14648
rect 10782 12960 10838 13016
rect 10874 12844 10930 12880
rect 10874 12824 10876 12844
rect 10876 12824 10928 12844
rect 10928 12824 10930 12844
rect 11058 12824 11114 12880
rect 10598 12416 10654 12472
rect 10046 8608 10102 8664
rect 9954 8064 10010 8120
rect 9862 6568 9918 6624
rect 9678 4528 9734 4584
rect 8850 2760 8906 2816
rect 9034 2644 9090 2680
rect 9034 2624 9036 2644
rect 9036 2624 9088 2644
rect 9088 2624 9090 2644
rect 8482 2352 8538 2408
rect 9678 4120 9734 4176
rect 9586 4020 9588 4040
rect 9588 4020 9640 4040
rect 9640 4020 9642 4040
rect 9586 3984 9642 4020
rect 9494 3168 9550 3224
rect 9954 6432 10010 6488
rect 10874 11772 10876 11792
rect 10876 11772 10928 11792
rect 10928 11772 10930 11792
rect 10874 11736 10930 11772
rect 12616 17434 12672 17436
rect 12696 17434 12752 17436
rect 12776 17434 12832 17436
rect 12856 17434 12912 17436
rect 12616 17382 12662 17434
rect 12662 17382 12672 17434
rect 12696 17382 12726 17434
rect 12726 17382 12738 17434
rect 12738 17382 12752 17434
rect 12776 17382 12790 17434
rect 12790 17382 12802 17434
rect 12802 17382 12832 17434
rect 12856 17382 12866 17434
rect 12866 17382 12912 17434
rect 12616 17380 12672 17382
rect 12696 17380 12752 17382
rect 12776 17380 12832 17382
rect 12856 17380 12912 17382
rect 12438 17312 12494 17368
rect 12346 16904 12402 16960
rect 11956 16890 12012 16892
rect 12036 16890 12092 16892
rect 12116 16890 12172 16892
rect 12196 16890 12252 16892
rect 11956 16838 12002 16890
rect 12002 16838 12012 16890
rect 12036 16838 12066 16890
rect 12066 16838 12078 16890
rect 12078 16838 12092 16890
rect 12116 16838 12130 16890
rect 12130 16838 12142 16890
rect 12142 16838 12172 16890
rect 12196 16838 12206 16890
rect 12206 16838 12252 16890
rect 11956 16836 12012 16838
rect 12036 16836 12092 16838
rect 12116 16836 12172 16838
rect 12196 16836 12252 16838
rect 12438 16768 12494 16824
rect 11794 16360 11850 16416
rect 12616 16346 12672 16348
rect 12696 16346 12752 16348
rect 12776 16346 12832 16348
rect 12856 16346 12912 16348
rect 12616 16294 12662 16346
rect 12662 16294 12672 16346
rect 12696 16294 12726 16346
rect 12726 16294 12738 16346
rect 12738 16294 12752 16346
rect 12776 16294 12790 16346
rect 12790 16294 12802 16346
rect 12802 16294 12832 16346
rect 12856 16294 12866 16346
rect 12866 16294 12912 16346
rect 12616 16292 12672 16294
rect 12696 16292 12752 16294
rect 12776 16292 12832 16294
rect 12856 16292 12912 16294
rect 12254 16088 12310 16144
rect 11426 15136 11482 15192
rect 11518 14456 11574 14512
rect 11426 13776 11482 13832
rect 11242 13268 11244 13288
rect 11244 13268 11296 13288
rect 11296 13268 11298 13288
rect 11242 13232 11298 13268
rect 11242 12960 11298 13016
rect 11334 12688 11390 12744
rect 10966 11328 11022 11384
rect 10966 11192 11022 11248
rect 10966 10784 11022 10840
rect 10966 10648 11022 10704
rect 10506 9016 10562 9072
rect 10414 8472 10470 8528
rect 9862 2896 9918 2952
rect 8390 1128 8446 1184
rect 7378 992 7434 1048
rect 11058 9832 11114 9888
rect 10782 9152 10838 9208
rect 10782 8472 10838 8528
rect 10966 9016 11022 9072
rect 10782 6976 10838 7032
rect 11956 15802 12012 15804
rect 12036 15802 12092 15804
rect 12116 15802 12172 15804
rect 12196 15802 12252 15804
rect 11956 15750 12002 15802
rect 12002 15750 12012 15802
rect 12036 15750 12066 15802
rect 12066 15750 12078 15802
rect 12078 15750 12092 15802
rect 12116 15750 12130 15802
rect 12130 15750 12142 15802
rect 12142 15750 12172 15802
rect 12196 15750 12206 15802
rect 12206 15750 12252 15802
rect 11956 15748 12012 15750
rect 12036 15748 12092 15750
rect 12116 15748 12172 15750
rect 12196 15748 12252 15750
rect 12346 15680 12402 15736
rect 11702 15136 11758 15192
rect 11702 13504 11758 13560
rect 11956 14714 12012 14716
rect 12036 14714 12092 14716
rect 12116 14714 12172 14716
rect 12196 14714 12252 14716
rect 11956 14662 12002 14714
rect 12002 14662 12012 14714
rect 12036 14662 12066 14714
rect 12066 14662 12078 14714
rect 12078 14662 12092 14714
rect 12116 14662 12130 14714
rect 12130 14662 12142 14714
rect 12142 14662 12172 14714
rect 12196 14662 12206 14714
rect 12206 14662 12252 14714
rect 11956 14660 12012 14662
rect 12036 14660 12092 14662
rect 12116 14660 12172 14662
rect 12196 14660 12252 14662
rect 12070 14456 12126 14512
rect 12070 14184 12126 14240
rect 11886 13912 11942 13968
rect 11956 13626 12012 13628
rect 12036 13626 12092 13628
rect 12116 13626 12172 13628
rect 12196 13626 12252 13628
rect 11956 13574 12002 13626
rect 12002 13574 12012 13626
rect 12036 13574 12066 13626
rect 12066 13574 12078 13626
rect 12078 13574 12092 13626
rect 12116 13574 12130 13626
rect 12130 13574 12142 13626
rect 12142 13574 12172 13626
rect 12196 13574 12206 13626
rect 12206 13574 12252 13626
rect 11956 13572 12012 13574
rect 12036 13572 12092 13574
rect 12116 13572 12172 13574
rect 12196 13572 12252 13574
rect 12438 14048 12494 14104
rect 12806 15444 12808 15464
rect 12808 15444 12860 15464
rect 12860 15444 12862 15464
rect 12806 15408 12862 15444
rect 12616 15258 12672 15260
rect 12696 15258 12752 15260
rect 12776 15258 12832 15260
rect 12856 15258 12912 15260
rect 12616 15206 12662 15258
rect 12662 15206 12672 15258
rect 12696 15206 12726 15258
rect 12726 15206 12738 15258
rect 12738 15206 12752 15258
rect 12776 15206 12790 15258
rect 12790 15206 12802 15258
rect 12802 15206 12832 15258
rect 12856 15206 12866 15258
rect 12866 15206 12912 15258
rect 12616 15204 12672 15206
rect 12696 15204 12752 15206
rect 12776 15204 12832 15206
rect 12856 15204 12912 15206
rect 12806 14592 12862 14648
rect 12990 14728 13046 14784
rect 12616 14170 12672 14172
rect 12696 14170 12752 14172
rect 12776 14170 12832 14172
rect 12856 14170 12912 14172
rect 12616 14118 12662 14170
rect 12662 14118 12672 14170
rect 12696 14118 12726 14170
rect 12726 14118 12738 14170
rect 12738 14118 12752 14170
rect 12776 14118 12790 14170
rect 12790 14118 12802 14170
rect 12802 14118 12832 14170
rect 12856 14118 12866 14170
rect 12866 14118 12912 14170
rect 12616 14116 12672 14118
rect 12696 14116 12752 14118
rect 12776 14116 12832 14118
rect 12856 14116 12912 14118
rect 11702 12824 11758 12880
rect 11610 12688 11666 12744
rect 11518 12552 11574 12608
rect 11242 10512 11298 10568
rect 11956 12538 12012 12540
rect 12036 12538 12092 12540
rect 12116 12538 12172 12540
rect 12196 12538 12252 12540
rect 11956 12486 12002 12538
rect 12002 12486 12012 12538
rect 12036 12486 12066 12538
rect 12066 12486 12078 12538
rect 12078 12486 12092 12538
rect 12116 12486 12130 12538
rect 12130 12486 12142 12538
rect 12142 12486 12172 12538
rect 12196 12486 12206 12538
rect 12206 12486 12252 12538
rect 11956 12484 12012 12486
rect 12036 12484 12092 12486
rect 12116 12484 12172 12486
rect 12196 12484 12252 12486
rect 11794 12416 11850 12472
rect 11794 11736 11850 11792
rect 12438 11872 12494 11928
rect 11956 11450 12012 11452
rect 12036 11450 12092 11452
rect 12116 11450 12172 11452
rect 12196 11450 12252 11452
rect 11956 11398 12002 11450
rect 12002 11398 12012 11450
rect 12036 11398 12066 11450
rect 12066 11398 12078 11450
rect 12078 11398 12092 11450
rect 12116 11398 12130 11450
rect 12130 11398 12142 11450
rect 12142 11398 12172 11450
rect 12196 11398 12206 11450
rect 12206 11398 12252 11450
rect 11956 11396 12012 11398
rect 12036 11396 12092 11398
rect 12116 11396 12172 11398
rect 12196 11396 12252 11398
rect 11058 6976 11114 7032
rect 10874 5480 10930 5536
rect 10782 4936 10838 4992
rect 10966 3984 11022 4040
rect 10782 2896 10838 2952
rect 11334 7928 11390 7984
rect 11518 10668 11574 10704
rect 11518 10648 11520 10668
rect 11520 10648 11572 10668
rect 11572 10648 11574 10668
rect 12070 11056 12126 11112
rect 12438 11328 12494 11384
rect 12616 13082 12672 13084
rect 12696 13082 12752 13084
rect 12776 13082 12832 13084
rect 12856 13082 12912 13084
rect 12616 13030 12662 13082
rect 12662 13030 12672 13082
rect 12696 13030 12726 13082
rect 12726 13030 12738 13082
rect 12738 13030 12752 13082
rect 12776 13030 12790 13082
rect 12790 13030 12802 13082
rect 12802 13030 12832 13082
rect 12856 13030 12866 13082
rect 12866 13030 12912 13082
rect 12616 13028 12672 13030
rect 12696 13028 12752 13030
rect 12776 13028 12832 13030
rect 12856 13028 12912 13030
rect 13174 14048 13230 14104
rect 13082 12960 13138 13016
rect 13910 16904 13966 16960
rect 13358 14864 13414 14920
rect 12990 12180 12992 12200
rect 12992 12180 13044 12200
rect 13044 12180 13046 12200
rect 12990 12144 13046 12180
rect 12616 11994 12672 11996
rect 12696 11994 12752 11996
rect 12776 11994 12832 11996
rect 12856 11994 12912 11996
rect 12616 11942 12662 11994
rect 12662 11942 12672 11994
rect 12696 11942 12726 11994
rect 12726 11942 12738 11994
rect 12738 11942 12752 11994
rect 12776 11942 12790 11994
rect 12790 11942 12802 11994
rect 12802 11942 12832 11994
rect 12856 11942 12866 11994
rect 12866 11942 12912 11994
rect 12616 11940 12672 11942
rect 12696 11940 12752 11942
rect 12776 11940 12832 11942
rect 12856 11940 12912 11942
rect 12616 10906 12672 10908
rect 12696 10906 12752 10908
rect 12776 10906 12832 10908
rect 12856 10906 12912 10908
rect 12616 10854 12662 10906
rect 12662 10854 12672 10906
rect 12696 10854 12726 10906
rect 12726 10854 12738 10906
rect 12738 10854 12752 10906
rect 12776 10854 12790 10906
rect 12790 10854 12802 10906
rect 12802 10854 12832 10906
rect 12856 10854 12866 10906
rect 12866 10854 12912 10906
rect 12616 10852 12672 10854
rect 12696 10852 12752 10854
rect 12776 10852 12832 10854
rect 12856 10852 12912 10854
rect 12438 10784 12494 10840
rect 11956 10362 12012 10364
rect 12036 10362 12092 10364
rect 12116 10362 12172 10364
rect 12196 10362 12252 10364
rect 11956 10310 12002 10362
rect 12002 10310 12012 10362
rect 12036 10310 12066 10362
rect 12066 10310 12078 10362
rect 12078 10310 12092 10362
rect 12116 10310 12130 10362
rect 12130 10310 12142 10362
rect 12142 10310 12172 10362
rect 12196 10310 12206 10362
rect 12206 10310 12252 10362
rect 11956 10308 12012 10310
rect 12036 10308 12092 10310
rect 12116 10308 12172 10310
rect 12196 10308 12252 10310
rect 11794 10240 11850 10296
rect 11610 9036 11666 9072
rect 11610 9016 11612 9036
rect 11612 9016 11664 9036
rect 11664 9016 11666 9036
rect 11610 7656 11666 7712
rect 11610 7112 11666 7168
rect 12254 9968 12310 10024
rect 12162 9716 12218 9752
rect 12162 9696 12164 9716
rect 12164 9696 12216 9716
rect 12216 9696 12218 9716
rect 11956 9274 12012 9276
rect 12036 9274 12092 9276
rect 12116 9274 12172 9276
rect 12196 9274 12252 9276
rect 11956 9222 12002 9274
rect 12002 9222 12012 9274
rect 12036 9222 12066 9274
rect 12066 9222 12078 9274
rect 12078 9222 12092 9274
rect 12116 9222 12130 9274
rect 12130 9222 12142 9274
rect 12142 9222 12172 9274
rect 12196 9222 12206 9274
rect 12206 9222 12252 9274
rect 11956 9220 12012 9222
rect 12036 9220 12092 9222
rect 12116 9220 12172 9222
rect 12196 9220 12252 9222
rect 11886 8472 11942 8528
rect 12254 8744 12310 8800
rect 11956 8186 12012 8188
rect 12036 8186 12092 8188
rect 12116 8186 12172 8188
rect 12196 8186 12252 8188
rect 11956 8134 12002 8186
rect 12002 8134 12012 8186
rect 12036 8134 12066 8186
rect 12066 8134 12078 8186
rect 12078 8134 12092 8186
rect 12116 8134 12130 8186
rect 12130 8134 12142 8186
rect 12142 8134 12172 8186
rect 12196 8134 12206 8186
rect 12206 8134 12252 8186
rect 11956 8132 12012 8134
rect 12036 8132 12092 8134
rect 12116 8132 12172 8134
rect 12196 8132 12252 8134
rect 12714 10376 12770 10432
rect 13174 12180 13176 12200
rect 13176 12180 13228 12200
rect 13228 12180 13230 12200
rect 13174 12144 13230 12180
rect 13450 13776 13506 13832
rect 13266 11464 13322 11520
rect 12616 9818 12672 9820
rect 12696 9818 12752 9820
rect 12776 9818 12832 9820
rect 12856 9818 12912 9820
rect 12616 9766 12662 9818
rect 12662 9766 12672 9818
rect 12696 9766 12726 9818
rect 12726 9766 12738 9818
rect 12738 9766 12752 9818
rect 12776 9766 12790 9818
rect 12790 9766 12802 9818
rect 12802 9766 12832 9818
rect 12856 9766 12866 9818
rect 12866 9766 12912 9818
rect 12616 9764 12672 9766
rect 12696 9764 12752 9766
rect 12776 9764 12832 9766
rect 12856 9764 12912 9766
rect 12530 9016 12586 9072
rect 11978 7404 12034 7440
rect 11978 7384 11980 7404
rect 11980 7384 12032 7404
rect 12032 7384 12034 7404
rect 11956 7098 12012 7100
rect 12036 7098 12092 7100
rect 12116 7098 12172 7100
rect 12196 7098 12252 7100
rect 11956 7046 12002 7098
rect 12002 7046 12012 7098
rect 12036 7046 12066 7098
rect 12066 7046 12078 7098
rect 12078 7046 12092 7098
rect 12116 7046 12130 7098
rect 12130 7046 12142 7098
rect 12142 7046 12172 7098
rect 12196 7046 12206 7098
rect 12206 7046 12252 7098
rect 11956 7044 12012 7046
rect 12036 7044 12092 7046
rect 12116 7044 12172 7046
rect 12196 7044 12252 7046
rect 11956 6010 12012 6012
rect 12036 6010 12092 6012
rect 12116 6010 12172 6012
rect 12196 6010 12252 6012
rect 11956 5958 12002 6010
rect 12002 5958 12012 6010
rect 12036 5958 12066 6010
rect 12066 5958 12078 6010
rect 12078 5958 12092 6010
rect 12116 5958 12130 6010
rect 12130 5958 12142 6010
rect 12142 5958 12172 6010
rect 12196 5958 12206 6010
rect 12206 5958 12252 6010
rect 11956 5956 12012 5958
rect 12036 5956 12092 5958
rect 12116 5956 12172 5958
rect 12196 5956 12252 5958
rect 11518 5208 11574 5264
rect 11794 5480 11850 5536
rect 12254 5344 12310 5400
rect 11956 4922 12012 4924
rect 12036 4922 12092 4924
rect 12116 4922 12172 4924
rect 12196 4922 12252 4924
rect 11956 4870 12002 4922
rect 12002 4870 12012 4922
rect 12036 4870 12066 4922
rect 12066 4870 12078 4922
rect 12078 4870 12092 4922
rect 12116 4870 12130 4922
rect 12130 4870 12142 4922
rect 12142 4870 12172 4922
rect 12196 4870 12206 4922
rect 12206 4870 12252 4922
rect 11956 4868 12012 4870
rect 12036 4868 12092 4870
rect 12116 4868 12172 4870
rect 12196 4868 12252 4870
rect 12616 8730 12672 8732
rect 12696 8730 12752 8732
rect 12776 8730 12832 8732
rect 12856 8730 12912 8732
rect 12616 8678 12662 8730
rect 12662 8678 12672 8730
rect 12696 8678 12726 8730
rect 12726 8678 12738 8730
rect 12738 8678 12752 8730
rect 12776 8678 12790 8730
rect 12790 8678 12802 8730
rect 12802 8678 12832 8730
rect 12856 8678 12866 8730
rect 12866 8678 12912 8730
rect 12616 8676 12672 8678
rect 12696 8676 12752 8678
rect 12776 8676 12832 8678
rect 12856 8676 12912 8678
rect 12622 8064 12678 8120
rect 12990 8200 13046 8256
rect 12616 7642 12672 7644
rect 12696 7642 12752 7644
rect 12776 7642 12832 7644
rect 12856 7642 12912 7644
rect 12616 7590 12662 7642
rect 12662 7590 12672 7642
rect 12696 7590 12726 7642
rect 12726 7590 12738 7642
rect 12738 7590 12752 7642
rect 12776 7590 12790 7642
rect 12790 7590 12802 7642
rect 12802 7590 12832 7642
rect 12856 7590 12866 7642
rect 12866 7590 12912 7642
rect 12616 7588 12672 7590
rect 12696 7588 12752 7590
rect 12776 7588 12832 7590
rect 12856 7588 12912 7590
rect 13266 10804 13322 10840
rect 13266 10784 13268 10804
rect 13268 10784 13320 10804
rect 13320 10784 13322 10804
rect 13266 9716 13322 9752
rect 13266 9696 13268 9716
rect 13268 9696 13320 9716
rect 13320 9696 13322 9716
rect 12622 6840 12678 6896
rect 12616 6554 12672 6556
rect 12696 6554 12752 6556
rect 12776 6554 12832 6556
rect 12856 6554 12912 6556
rect 12616 6502 12662 6554
rect 12662 6502 12672 6554
rect 12696 6502 12726 6554
rect 12726 6502 12738 6554
rect 12738 6502 12752 6554
rect 12776 6502 12790 6554
rect 12790 6502 12802 6554
rect 12802 6502 12832 6554
rect 12856 6502 12866 6554
rect 12866 6502 12912 6554
rect 12616 6500 12672 6502
rect 12696 6500 12752 6502
rect 12776 6500 12832 6502
rect 12856 6500 12912 6502
rect 12438 5888 12494 5944
rect 12714 6024 12770 6080
rect 12616 5466 12672 5468
rect 12696 5466 12752 5468
rect 12776 5466 12832 5468
rect 12856 5466 12912 5468
rect 12616 5414 12662 5466
rect 12662 5414 12672 5466
rect 12696 5414 12726 5466
rect 12726 5414 12738 5466
rect 12738 5414 12752 5466
rect 12776 5414 12790 5466
rect 12790 5414 12802 5466
rect 12802 5414 12832 5466
rect 12856 5414 12866 5466
rect 12866 5414 12912 5466
rect 12616 5412 12672 5414
rect 12696 5412 12752 5414
rect 12776 5412 12832 5414
rect 12856 5412 12912 5414
rect 12438 4800 12494 4856
rect 11794 4564 11796 4584
rect 11796 4564 11848 4584
rect 11848 4564 11850 4584
rect 11794 4528 11850 4564
rect 12438 4392 12494 4448
rect 12990 4528 13046 4584
rect 12616 4378 12672 4380
rect 12696 4378 12752 4380
rect 12776 4378 12832 4380
rect 12856 4378 12912 4380
rect 12616 4326 12662 4378
rect 12662 4326 12672 4378
rect 12696 4326 12726 4378
rect 12726 4326 12738 4378
rect 12738 4326 12752 4378
rect 12776 4326 12790 4378
rect 12790 4326 12802 4378
rect 12802 4326 12832 4378
rect 12856 4326 12866 4378
rect 12866 4326 12912 4378
rect 12616 4324 12672 4326
rect 12696 4324 12752 4326
rect 12776 4324 12832 4326
rect 12856 4324 12912 4326
rect 12346 4140 12402 4176
rect 12346 4120 12348 4140
rect 12348 4120 12400 4140
rect 12400 4120 12402 4140
rect 10322 1672 10378 1728
rect 11334 2388 11336 2408
rect 11336 2388 11388 2408
rect 11388 2388 11390 2408
rect 11334 2352 11390 2388
rect 11702 3848 11758 3904
rect 11702 3576 11758 3632
rect 11956 3834 12012 3836
rect 12036 3834 12092 3836
rect 12116 3834 12172 3836
rect 12196 3834 12252 3836
rect 11956 3782 12002 3834
rect 12002 3782 12012 3834
rect 12036 3782 12066 3834
rect 12066 3782 12078 3834
rect 12078 3782 12092 3834
rect 12116 3782 12130 3834
rect 12130 3782 12142 3834
rect 12142 3782 12172 3834
rect 12196 3782 12206 3834
rect 12206 3782 12252 3834
rect 11956 3780 12012 3782
rect 12036 3780 12092 3782
rect 12116 3780 12172 3782
rect 12196 3780 12252 3782
rect 12346 3712 12402 3768
rect 3882 448 3938 504
rect 12806 3612 12808 3632
rect 12808 3612 12860 3632
rect 12860 3612 12862 3632
rect 12806 3576 12862 3612
rect 12346 3304 12402 3360
rect 12438 3168 12494 3224
rect 11956 2746 12012 2748
rect 12036 2746 12092 2748
rect 12116 2746 12172 2748
rect 12196 2746 12252 2748
rect 11956 2694 12002 2746
rect 12002 2694 12012 2746
rect 12036 2694 12066 2746
rect 12066 2694 12078 2746
rect 12078 2694 12092 2746
rect 12116 2694 12130 2746
rect 12130 2694 12142 2746
rect 12142 2694 12172 2746
rect 12196 2694 12206 2746
rect 12206 2694 12252 2746
rect 11956 2692 12012 2694
rect 12036 2692 12092 2694
rect 12116 2692 12172 2694
rect 12196 2692 12252 2694
rect 11978 2488 12034 2544
rect 12346 720 12402 776
rect 12616 3290 12672 3292
rect 12696 3290 12752 3292
rect 12776 3290 12832 3292
rect 12856 3290 12912 3292
rect 12616 3238 12662 3290
rect 12662 3238 12672 3290
rect 12696 3238 12726 3290
rect 12726 3238 12738 3290
rect 12738 3238 12752 3290
rect 12776 3238 12790 3290
rect 12790 3238 12802 3290
rect 12802 3238 12832 3290
rect 12856 3238 12866 3290
rect 12866 3238 12912 3290
rect 12616 3236 12672 3238
rect 12696 3236 12752 3238
rect 12776 3236 12832 3238
rect 12856 3236 12912 3238
rect 13450 7112 13506 7168
rect 14002 11872 14058 11928
rect 13910 11464 13966 11520
rect 13910 11328 13966 11384
rect 13818 11056 13874 11112
rect 13726 8200 13782 8256
rect 13910 7928 13966 7984
rect 13634 6568 13690 6624
rect 13634 4800 13690 4856
rect 13542 4392 13598 4448
rect 12616 2202 12672 2204
rect 12696 2202 12752 2204
rect 12776 2202 12832 2204
rect 12856 2202 12912 2204
rect 12616 2150 12662 2202
rect 12662 2150 12672 2202
rect 12696 2150 12726 2202
rect 12726 2150 12738 2202
rect 12738 2150 12752 2202
rect 12776 2150 12790 2202
rect 12790 2150 12802 2202
rect 12802 2150 12832 2202
rect 12856 2150 12866 2202
rect 12866 2150 12912 2202
rect 12616 2148 12672 2150
rect 12696 2148 12752 2150
rect 12776 2148 12832 2150
rect 12856 2148 12912 2150
rect 13726 2624 13782 2680
rect 14278 14456 14334 14512
rect 14186 13368 14242 13424
rect 14554 16632 14610 16688
rect 14278 12280 14334 12336
rect 14186 12144 14242 12200
rect 14278 12008 14334 12064
rect 14186 11348 14242 11384
rect 14186 11328 14188 11348
rect 14188 11328 14240 11348
rect 14240 11328 14242 11348
rect 14186 10104 14242 10160
rect 14186 9832 14242 9888
rect 14370 11464 14426 11520
rect 14278 9324 14280 9344
rect 14280 9324 14332 9344
rect 14332 9324 14334 9344
rect 14278 9288 14334 9324
rect 14186 5616 14242 5672
rect 15198 16496 15254 16552
rect 14830 15680 14886 15736
rect 14738 13776 14794 13832
rect 14554 12280 14610 12336
rect 14554 10784 14610 10840
rect 14462 10240 14518 10296
rect 14554 10104 14610 10160
rect 14462 9288 14518 9344
rect 14554 8472 14610 8528
rect 14370 7112 14426 7168
rect 14830 11464 14886 11520
rect 14830 10784 14886 10840
rect 14922 8744 14978 8800
rect 14830 7656 14886 7712
rect 14738 7112 14794 7168
rect 14554 5072 14610 5128
rect 14646 4664 14702 4720
rect 14830 4800 14886 4856
rect 11610 584 11666 640
rect 15474 13268 15476 13288
rect 15476 13268 15528 13288
rect 15528 13268 15530 13288
rect 15474 13232 15530 13268
rect 15290 10784 15346 10840
rect 15198 10240 15254 10296
rect 17498 18536 17554 18592
rect 17406 18400 17462 18456
rect 15658 12552 15714 12608
rect 15106 9580 15162 9616
rect 15106 9560 15108 9580
rect 15108 9560 15160 9580
rect 15160 9560 15162 9580
rect 15106 8064 15162 8120
rect 15566 9424 15622 9480
rect 15382 6976 15438 7032
rect 15382 6704 15438 6760
rect 15382 3032 15438 3088
rect 15290 992 15346 1048
rect 15658 8880 15714 8936
rect 15934 12552 15990 12608
rect 16394 15000 16450 15056
rect 17314 17196 17370 17232
rect 17314 17176 17316 17196
rect 17316 17176 17368 17196
rect 17368 17176 17370 17196
rect 16956 16890 17012 16892
rect 17036 16890 17092 16892
rect 17116 16890 17172 16892
rect 17196 16890 17252 16892
rect 16956 16838 17002 16890
rect 17002 16838 17012 16890
rect 17036 16838 17066 16890
rect 17066 16838 17078 16890
rect 17078 16838 17092 16890
rect 17116 16838 17130 16890
rect 17130 16838 17142 16890
rect 17142 16838 17172 16890
rect 17196 16838 17206 16890
rect 17206 16838 17252 16890
rect 16956 16836 17012 16838
rect 17036 16836 17092 16838
rect 17116 16836 17172 16838
rect 17196 16836 17252 16838
rect 17130 16532 17132 16552
rect 17132 16532 17184 16552
rect 17184 16532 17186 16552
rect 16302 12960 16358 13016
rect 17130 16496 17186 16532
rect 17038 16088 17094 16144
rect 16956 15802 17012 15804
rect 17036 15802 17092 15804
rect 17116 15802 17172 15804
rect 17196 15802 17252 15804
rect 16956 15750 17002 15802
rect 17002 15750 17012 15802
rect 17036 15750 17066 15802
rect 17066 15750 17078 15802
rect 17078 15750 17092 15802
rect 17116 15750 17130 15802
rect 17130 15750 17142 15802
rect 17142 15750 17172 15802
rect 17196 15750 17206 15802
rect 17206 15750 17252 15802
rect 16956 15748 17012 15750
rect 17036 15748 17092 15750
rect 17116 15748 17172 15750
rect 17196 15748 17252 15750
rect 16956 14714 17012 14716
rect 17036 14714 17092 14716
rect 17116 14714 17172 14716
rect 17196 14714 17252 14716
rect 16956 14662 17002 14714
rect 17002 14662 17012 14714
rect 17036 14662 17066 14714
rect 17066 14662 17078 14714
rect 17078 14662 17092 14714
rect 17116 14662 17130 14714
rect 17130 14662 17142 14714
rect 17142 14662 17172 14714
rect 17196 14662 17206 14714
rect 17206 14662 17252 14714
rect 16956 14660 17012 14662
rect 17036 14660 17092 14662
rect 17116 14660 17172 14662
rect 17196 14660 17252 14662
rect 16956 13626 17012 13628
rect 17036 13626 17092 13628
rect 17116 13626 17172 13628
rect 17196 13626 17252 13628
rect 16956 13574 17002 13626
rect 17002 13574 17012 13626
rect 17036 13574 17066 13626
rect 17066 13574 17078 13626
rect 17078 13574 17092 13626
rect 17116 13574 17130 13626
rect 17130 13574 17142 13626
rect 17142 13574 17172 13626
rect 17196 13574 17206 13626
rect 17206 13574 17252 13626
rect 16956 13572 17012 13574
rect 17036 13572 17092 13574
rect 17116 13572 17172 13574
rect 17196 13572 17252 13574
rect 15842 11228 15844 11248
rect 15844 11228 15896 11248
rect 15896 11228 15898 11248
rect 15842 11192 15898 11228
rect 15934 10784 15990 10840
rect 15934 10376 15990 10432
rect 15842 10240 15898 10296
rect 16210 7948 16266 7984
rect 16210 7928 16212 7948
rect 16212 7928 16264 7948
rect 16264 7928 16266 7948
rect 16486 12180 16488 12200
rect 16488 12180 16540 12200
rect 16540 12180 16542 12200
rect 16486 12144 16542 12180
rect 16486 9696 16542 9752
rect 16670 11736 16726 11792
rect 16956 12538 17012 12540
rect 17036 12538 17092 12540
rect 17116 12538 17172 12540
rect 17196 12538 17252 12540
rect 16956 12486 17002 12538
rect 17002 12486 17012 12538
rect 17036 12486 17066 12538
rect 17066 12486 17078 12538
rect 17078 12486 17092 12538
rect 17116 12486 17130 12538
rect 17130 12486 17142 12538
rect 17142 12486 17172 12538
rect 17196 12486 17206 12538
rect 17206 12486 17252 12538
rect 16956 12484 17012 12486
rect 17036 12484 17092 12486
rect 17116 12484 17172 12486
rect 17196 12484 17252 12486
rect 16956 11450 17012 11452
rect 17036 11450 17092 11452
rect 17116 11450 17172 11452
rect 17196 11450 17252 11452
rect 16956 11398 17002 11450
rect 17002 11398 17012 11450
rect 17036 11398 17066 11450
rect 17066 11398 17078 11450
rect 17078 11398 17092 11450
rect 17116 11398 17130 11450
rect 17130 11398 17142 11450
rect 17142 11398 17172 11450
rect 17196 11398 17206 11450
rect 17206 11398 17252 11450
rect 16956 11396 17012 11398
rect 17036 11396 17092 11398
rect 17116 11396 17172 11398
rect 17196 11396 17252 11398
rect 17038 10920 17094 10976
rect 16762 10104 16818 10160
rect 16486 9580 16542 9616
rect 16486 9560 16488 9580
rect 16488 9560 16540 9580
rect 16540 9560 16542 9580
rect 15658 4120 15714 4176
rect 16026 6296 16082 6352
rect 15934 5480 15990 5536
rect 15934 4392 15990 4448
rect 16210 6568 16266 6624
rect 16210 6432 16266 6488
rect 16026 4120 16082 4176
rect 15566 2896 15622 2952
rect 16118 3304 16174 3360
rect 16486 6024 16542 6080
rect 16578 5888 16634 5944
rect 16302 4392 16358 4448
rect 16956 10362 17012 10364
rect 17036 10362 17092 10364
rect 17116 10362 17172 10364
rect 17196 10362 17252 10364
rect 16956 10310 17002 10362
rect 17002 10310 17012 10362
rect 17036 10310 17066 10362
rect 17066 10310 17078 10362
rect 17078 10310 17092 10362
rect 17116 10310 17130 10362
rect 17130 10310 17142 10362
rect 17142 10310 17172 10362
rect 17196 10310 17206 10362
rect 17206 10310 17252 10362
rect 16956 10308 17012 10310
rect 17036 10308 17092 10310
rect 17116 10308 17172 10310
rect 17196 10308 17252 10310
rect 17038 9832 17094 9888
rect 16956 9274 17012 9276
rect 17036 9274 17092 9276
rect 17116 9274 17172 9276
rect 17196 9274 17252 9276
rect 16956 9222 17002 9274
rect 17002 9222 17012 9274
rect 17036 9222 17066 9274
rect 17066 9222 17078 9274
rect 17078 9222 17092 9274
rect 17116 9222 17130 9274
rect 17130 9222 17142 9274
rect 17142 9222 17172 9274
rect 17196 9222 17206 9274
rect 17206 9222 17252 9274
rect 16956 9220 17012 9222
rect 17036 9220 17092 9222
rect 17116 9220 17172 9222
rect 17196 9220 17252 9222
rect 16956 8186 17012 8188
rect 17036 8186 17092 8188
rect 17116 8186 17172 8188
rect 17196 8186 17252 8188
rect 16956 8134 17002 8186
rect 17002 8134 17012 8186
rect 17036 8134 17066 8186
rect 17066 8134 17078 8186
rect 17078 8134 17092 8186
rect 17116 8134 17130 8186
rect 17130 8134 17142 8186
rect 17142 8134 17172 8186
rect 17196 8134 17206 8186
rect 17206 8134 17252 8186
rect 16956 8132 17012 8134
rect 17036 8132 17092 8134
rect 17116 8132 17172 8134
rect 17196 8132 17252 8134
rect 17038 7828 17040 7848
rect 17040 7828 17092 7848
rect 17092 7828 17094 7848
rect 17038 7792 17094 7828
rect 17038 7248 17094 7304
rect 16956 7098 17012 7100
rect 17036 7098 17092 7100
rect 17116 7098 17172 7100
rect 17196 7098 17252 7100
rect 16956 7046 17002 7098
rect 17002 7046 17012 7098
rect 17036 7046 17066 7098
rect 17066 7046 17078 7098
rect 17078 7046 17092 7098
rect 17116 7046 17130 7098
rect 17130 7046 17142 7098
rect 17142 7046 17172 7098
rect 17196 7046 17206 7098
rect 17206 7046 17252 7098
rect 16956 7044 17012 7046
rect 17036 7044 17092 7046
rect 17116 7044 17172 7046
rect 17196 7044 17252 7046
rect 16762 6160 16818 6216
rect 16956 6010 17012 6012
rect 17036 6010 17092 6012
rect 17116 6010 17172 6012
rect 17196 6010 17252 6012
rect 16956 5958 17002 6010
rect 17002 5958 17012 6010
rect 17036 5958 17066 6010
rect 17066 5958 17078 6010
rect 17078 5958 17092 6010
rect 17116 5958 17130 6010
rect 17130 5958 17142 6010
rect 17142 5958 17172 6010
rect 17196 5958 17206 6010
rect 17206 5958 17252 6010
rect 16956 5956 17012 5958
rect 17036 5956 17092 5958
rect 17116 5956 17172 5958
rect 17196 5956 17252 5958
rect 18326 17720 18382 17776
rect 17616 17434 17672 17436
rect 17696 17434 17752 17436
rect 17776 17434 17832 17436
rect 17856 17434 17912 17436
rect 17616 17382 17662 17434
rect 17662 17382 17672 17434
rect 17696 17382 17726 17434
rect 17726 17382 17738 17434
rect 17738 17382 17752 17434
rect 17776 17382 17790 17434
rect 17790 17382 17802 17434
rect 17802 17382 17832 17434
rect 17856 17382 17866 17434
rect 17866 17382 17912 17434
rect 17616 17380 17672 17382
rect 17696 17380 17752 17382
rect 17776 17380 17832 17382
rect 17856 17380 17912 17382
rect 17616 16346 17672 16348
rect 17696 16346 17752 16348
rect 17776 16346 17832 16348
rect 17856 16346 17912 16348
rect 17616 16294 17662 16346
rect 17662 16294 17672 16346
rect 17696 16294 17726 16346
rect 17726 16294 17738 16346
rect 17738 16294 17752 16346
rect 17776 16294 17790 16346
rect 17790 16294 17802 16346
rect 17802 16294 17832 16346
rect 17856 16294 17866 16346
rect 17866 16294 17912 16346
rect 17616 16292 17672 16294
rect 17696 16292 17752 16294
rect 17776 16292 17832 16294
rect 17856 16292 17912 16294
rect 17616 15258 17672 15260
rect 17696 15258 17752 15260
rect 17776 15258 17832 15260
rect 17856 15258 17912 15260
rect 17616 15206 17662 15258
rect 17662 15206 17672 15258
rect 17696 15206 17726 15258
rect 17726 15206 17738 15258
rect 17738 15206 17752 15258
rect 17776 15206 17790 15258
rect 17790 15206 17802 15258
rect 17802 15206 17832 15258
rect 17856 15206 17866 15258
rect 17866 15206 17912 15258
rect 17616 15204 17672 15206
rect 17696 15204 17752 15206
rect 17776 15204 17832 15206
rect 17856 15204 17912 15206
rect 17616 14170 17672 14172
rect 17696 14170 17752 14172
rect 17776 14170 17832 14172
rect 17856 14170 17912 14172
rect 17616 14118 17662 14170
rect 17662 14118 17672 14170
rect 17696 14118 17726 14170
rect 17726 14118 17738 14170
rect 17738 14118 17752 14170
rect 17776 14118 17790 14170
rect 17790 14118 17802 14170
rect 17802 14118 17832 14170
rect 17856 14118 17866 14170
rect 17866 14118 17912 14170
rect 17616 14116 17672 14118
rect 17696 14116 17752 14118
rect 17776 14116 17832 14118
rect 17856 14116 17912 14118
rect 17498 13504 17554 13560
rect 17616 13082 17672 13084
rect 17696 13082 17752 13084
rect 17776 13082 17832 13084
rect 17856 13082 17912 13084
rect 17616 13030 17662 13082
rect 17662 13030 17672 13082
rect 17696 13030 17726 13082
rect 17726 13030 17738 13082
rect 17738 13030 17752 13082
rect 17776 13030 17790 13082
rect 17790 13030 17802 13082
rect 17802 13030 17832 13082
rect 17856 13030 17866 13082
rect 17866 13030 17912 13082
rect 17616 13028 17672 13030
rect 17696 13028 17752 13030
rect 17776 13028 17832 13030
rect 17856 13028 17912 13030
rect 17682 12844 17738 12880
rect 17682 12824 17684 12844
rect 17684 12824 17736 12844
rect 17736 12824 17738 12844
rect 17682 12688 17738 12744
rect 17406 11872 17462 11928
rect 18142 15544 18198 15600
rect 18418 16088 18474 16144
rect 18418 13640 18474 13696
rect 18234 12824 18290 12880
rect 17616 11994 17672 11996
rect 17696 11994 17752 11996
rect 17776 11994 17832 11996
rect 17856 11994 17912 11996
rect 17616 11942 17662 11994
rect 17662 11942 17672 11994
rect 17696 11942 17726 11994
rect 17726 11942 17738 11994
rect 17738 11942 17752 11994
rect 17776 11942 17790 11994
rect 17790 11942 17802 11994
rect 17802 11942 17832 11994
rect 17856 11942 17866 11994
rect 17866 11942 17912 11994
rect 17616 11940 17672 11942
rect 17696 11940 17752 11942
rect 17776 11940 17832 11942
rect 17856 11940 17912 11942
rect 17774 11192 17830 11248
rect 17958 11228 17960 11248
rect 17960 11228 18012 11248
rect 18012 11228 18014 11248
rect 17958 11192 18014 11228
rect 18326 11600 18382 11656
rect 18142 11056 18198 11112
rect 17616 10906 17672 10908
rect 17696 10906 17752 10908
rect 17776 10906 17832 10908
rect 17856 10906 17912 10908
rect 17616 10854 17662 10906
rect 17662 10854 17672 10906
rect 17696 10854 17726 10906
rect 17726 10854 17738 10906
rect 17738 10854 17752 10906
rect 17776 10854 17790 10906
rect 17790 10854 17802 10906
rect 17802 10854 17832 10906
rect 17856 10854 17866 10906
rect 17866 10854 17912 10906
rect 17616 10852 17672 10854
rect 17696 10852 17752 10854
rect 17776 10852 17832 10854
rect 17856 10852 17912 10854
rect 17958 10684 17960 10704
rect 17960 10684 18012 10704
rect 18012 10684 18014 10704
rect 17498 10532 17554 10568
rect 17498 10512 17500 10532
rect 17500 10512 17552 10532
rect 17552 10512 17554 10532
rect 17958 10648 18014 10684
rect 17774 10104 17830 10160
rect 17498 10004 17500 10024
rect 17500 10004 17552 10024
rect 17552 10004 17554 10024
rect 17498 9968 17554 10004
rect 17616 9818 17672 9820
rect 17696 9818 17752 9820
rect 17776 9818 17832 9820
rect 17856 9818 17912 9820
rect 17616 9766 17662 9818
rect 17662 9766 17672 9818
rect 17696 9766 17726 9818
rect 17726 9766 17738 9818
rect 17738 9766 17752 9818
rect 17776 9766 17790 9818
rect 17790 9766 17802 9818
rect 17802 9766 17832 9818
rect 17856 9766 17866 9818
rect 17866 9766 17912 9818
rect 17616 9764 17672 9766
rect 17696 9764 17752 9766
rect 17776 9764 17832 9766
rect 17856 9764 17912 9766
rect 16578 3304 16634 3360
rect 15842 856 15898 912
rect 16670 1672 16726 1728
rect 16956 4922 17012 4924
rect 17036 4922 17092 4924
rect 17116 4922 17172 4924
rect 17196 4922 17252 4924
rect 16956 4870 17002 4922
rect 17002 4870 17012 4922
rect 17036 4870 17066 4922
rect 17066 4870 17078 4922
rect 17078 4870 17092 4922
rect 17116 4870 17130 4922
rect 17130 4870 17142 4922
rect 17142 4870 17172 4922
rect 17196 4870 17206 4922
rect 17206 4870 17252 4922
rect 16956 4868 17012 4870
rect 17036 4868 17092 4870
rect 17116 4868 17172 4870
rect 17196 4868 17252 4870
rect 16956 3834 17012 3836
rect 17036 3834 17092 3836
rect 17116 3834 17172 3836
rect 17196 3834 17252 3836
rect 16956 3782 17002 3834
rect 17002 3782 17012 3834
rect 17036 3782 17066 3834
rect 17066 3782 17078 3834
rect 17078 3782 17092 3834
rect 17116 3782 17130 3834
rect 17130 3782 17142 3834
rect 17142 3782 17172 3834
rect 17196 3782 17206 3834
rect 17206 3782 17252 3834
rect 16956 3780 17012 3782
rect 17036 3780 17092 3782
rect 17116 3780 17172 3782
rect 17196 3780 17252 3782
rect 18142 10124 18198 10160
rect 18142 10104 18144 10124
rect 18144 10104 18196 10124
rect 18196 10104 18198 10124
rect 18142 9016 18198 9072
rect 18050 8880 18106 8936
rect 17616 8730 17672 8732
rect 17696 8730 17752 8732
rect 17776 8730 17832 8732
rect 17856 8730 17912 8732
rect 17616 8678 17662 8730
rect 17662 8678 17672 8730
rect 17696 8678 17726 8730
rect 17726 8678 17738 8730
rect 17738 8678 17752 8730
rect 17776 8678 17790 8730
rect 17790 8678 17802 8730
rect 17802 8678 17832 8730
rect 17856 8678 17866 8730
rect 17866 8678 17912 8730
rect 17616 8676 17672 8678
rect 17696 8676 17752 8678
rect 17776 8676 17832 8678
rect 17856 8676 17912 8678
rect 17590 7792 17646 7848
rect 17616 7642 17672 7644
rect 17696 7642 17752 7644
rect 17776 7642 17832 7644
rect 17856 7642 17912 7644
rect 17616 7590 17662 7642
rect 17662 7590 17672 7642
rect 17696 7590 17726 7642
rect 17726 7590 17738 7642
rect 17738 7590 17752 7642
rect 17776 7590 17790 7642
rect 17790 7590 17802 7642
rect 17802 7590 17832 7642
rect 17856 7590 17866 7642
rect 17866 7590 17912 7642
rect 17616 7588 17672 7590
rect 17696 7588 17752 7590
rect 17776 7588 17832 7590
rect 17856 7588 17912 7590
rect 17498 6840 17554 6896
rect 17616 6554 17672 6556
rect 17696 6554 17752 6556
rect 17776 6554 17832 6556
rect 17856 6554 17912 6556
rect 17616 6502 17662 6554
rect 17662 6502 17672 6554
rect 17696 6502 17726 6554
rect 17726 6502 17738 6554
rect 17738 6502 17752 6554
rect 17776 6502 17790 6554
rect 17790 6502 17802 6554
rect 17802 6502 17832 6554
rect 17856 6502 17866 6554
rect 17866 6502 17912 6554
rect 17616 6500 17672 6502
rect 17696 6500 17752 6502
rect 17776 6500 17832 6502
rect 17856 6500 17912 6502
rect 17616 5466 17672 5468
rect 17696 5466 17752 5468
rect 17776 5466 17832 5468
rect 17856 5466 17912 5468
rect 17616 5414 17662 5466
rect 17662 5414 17672 5466
rect 17696 5414 17726 5466
rect 17726 5414 17738 5466
rect 17738 5414 17752 5466
rect 17776 5414 17790 5466
rect 17790 5414 17802 5466
rect 17802 5414 17832 5466
rect 17856 5414 17866 5466
rect 17866 5414 17912 5466
rect 17616 5412 17672 5414
rect 17696 5412 17752 5414
rect 17776 5412 17832 5414
rect 17856 5412 17912 5414
rect 17616 4378 17672 4380
rect 17696 4378 17752 4380
rect 17776 4378 17832 4380
rect 17856 4378 17912 4380
rect 17616 4326 17662 4378
rect 17662 4326 17672 4378
rect 17696 4326 17726 4378
rect 17726 4326 17738 4378
rect 17738 4326 17752 4378
rect 17776 4326 17790 4378
rect 17790 4326 17802 4378
rect 17802 4326 17832 4378
rect 17856 4326 17866 4378
rect 17866 4326 17912 4378
rect 17616 4324 17672 4326
rect 17696 4324 17752 4326
rect 17776 4324 17832 4326
rect 17856 4324 17912 4326
rect 17958 3576 18014 3632
rect 18418 9696 18474 9752
rect 18418 8780 18420 8800
rect 18420 8780 18472 8800
rect 18472 8780 18474 8800
rect 18418 8744 18474 8780
rect 18418 6296 18474 6352
rect 18326 5480 18382 5536
rect 18234 3984 18290 4040
rect 16854 3304 16910 3360
rect 16956 2746 17012 2748
rect 17036 2746 17092 2748
rect 17116 2746 17172 2748
rect 17196 2746 17252 2748
rect 16956 2694 17002 2746
rect 17002 2694 17012 2746
rect 17036 2694 17066 2746
rect 17066 2694 17078 2746
rect 17078 2694 17092 2746
rect 17116 2694 17130 2746
rect 17130 2694 17142 2746
rect 17142 2694 17172 2746
rect 17196 2694 17206 2746
rect 17206 2694 17252 2746
rect 16956 2692 17012 2694
rect 17036 2692 17092 2694
rect 17116 2692 17172 2694
rect 17196 2692 17252 2694
rect 16946 2488 17002 2544
rect 17616 3290 17672 3292
rect 17696 3290 17752 3292
rect 17776 3290 17832 3292
rect 17856 3290 17912 3292
rect 17616 3238 17662 3290
rect 17662 3238 17672 3290
rect 17696 3238 17726 3290
rect 17726 3238 17738 3290
rect 17738 3238 17752 3290
rect 17776 3238 17790 3290
rect 17790 3238 17802 3290
rect 17802 3238 17832 3290
rect 17856 3238 17866 3290
rect 17866 3238 17912 3290
rect 17616 3236 17672 3238
rect 17696 3236 17752 3238
rect 17776 3236 17832 3238
rect 17856 3236 17912 3238
rect 18142 3476 18144 3496
rect 18144 3476 18196 3496
rect 18196 3476 18198 3496
rect 18142 3440 18198 3476
rect 18418 3884 18420 3904
rect 18420 3884 18472 3904
rect 18472 3884 18474 3904
rect 18418 3848 18474 3884
rect 18602 8472 18658 8528
rect 18878 8336 18934 8392
rect 19154 9424 19210 9480
rect 17958 2352 18014 2408
rect 17616 2202 17672 2204
rect 17696 2202 17752 2204
rect 17776 2202 17832 2204
rect 17856 2202 17912 2204
rect 17616 2150 17662 2202
rect 17662 2150 17672 2202
rect 17696 2150 17726 2202
rect 17726 2150 17738 2202
rect 17738 2150 17752 2202
rect 17776 2150 17790 2202
rect 17790 2150 17802 2202
rect 17802 2150 17832 2202
rect 17856 2150 17866 2202
rect 17866 2150 17912 2202
rect 17616 2148 17672 2150
rect 17696 2148 17752 2150
rect 17776 2148 17832 2150
rect 17856 2148 17912 2150
rect 18234 1536 18290 1592
rect 18326 1400 18382 1456
<< metal3 >>
rect 1117 18730 1183 18733
rect 15878 18730 15884 18732
rect 1117 18728 15884 18730
rect 1117 18672 1122 18728
rect 1178 18672 15884 18728
rect 1117 18670 15884 18672
rect 1117 18667 1183 18670
rect 15878 18668 15884 18670
rect 15948 18668 15954 18732
rect 0 18594 800 18624
rect 2957 18594 3023 18597
rect 0 18592 3023 18594
rect 0 18536 2962 18592
rect 3018 18536 3023 18592
rect 0 18534 3023 18536
rect 0 18504 800 18534
rect 2957 18531 3023 18534
rect 5022 18532 5028 18596
rect 5092 18594 5098 18596
rect 10869 18594 10935 18597
rect 5092 18592 10935 18594
rect 5092 18536 10874 18592
rect 10930 18536 10935 18592
rect 5092 18534 10935 18536
rect 5092 18532 5098 18534
rect 10869 18531 10935 18534
rect 17493 18594 17559 18597
rect 19200 18594 20000 18624
rect 17493 18592 20000 18594
rect 17493 18536 17498 18592
rect 17554 18536 20000 18592
rect 17493 18534 20000 18536
rect 17493 18531 17559 18534
rect 19200 18504 20000 18534
rect 1526 18396 1532 18460
rect 1596 18458 1602 18460
rect 17401 18458 17467 18461
rect 1596 18456 17467 18458
rect 1596 18400 17406 18456
rect 17462 18400 17467 18456
rect 1596 18398 17467 18400
rect 1596 18396 1602 18398
rect 17401 18395 17467 18398
rect 1301 18322 1367 18325
rect 13854 18322 13860 18324
rect 1301 18320 13860 18322
rect 1301 18264 1306 18320
rect 1362 18264 13860 18320
rect 1301 18262 13860 18264
rect 1301 18259 1367 18262
rect 13854 18260 13860 18262
rect 13924 18260 13930 18324
rect 6361 18186 6427 18189
rect 14590 18186 14596 18188
rect 6361 18184 14596 18186
rect 6361 18128 6366 18184
rect 6422 18128 14596 18184
rect 6361 18126 14596 18128
rect 6361 18123 6427 18126
rect 14590 18124 14596 18126
rect 14660 18124 14666 18188
rect 5809 18052 5875 18053
rect 5758 18050 5764 18052
rect 5718 17990 5764 18050
rect 5828 18048 5875 18052
rect 5870 17992 5875 18048
rect 5758 17988 5764 17990
rect 5828 17988 5875 17992
rect 5809 17987 5875 17988
rect 4245 17914 4311 17917
rect 12341 17914 12407 17917
rect 4245 17912 12407 17914
rect 4245 17856 4250 17912
rect 4306 17856 12346 17912
rect 12402 17856 12407 17912
rect 4245 17854 12407 17856
rect 4245 17851 4311 17854
rect 12341 17851 12407 17854
rect 749 17778 815 17781
rect 18321 17778 18387 17781
rect 749 17776 18387 17778
rect 749 17720 754 17776
rect 810 17720 18326 17776
rect 18382 17720 18387 17776
rect 749 17718 18387 17720
rect 749 17715 815 17718
rect 18321 17715 18387 17718
rect 2313 17642 2379 17645
rect 13486 17642 13492 17644
rect 2313 17640 13492 17642
rect 2313 17584 2318 17640
rect 2374 17584 13492 17640
rect 2313 17582 13492 17584
rect 2313 17579 2379 17582
rect 13486 17580 13492 17582
rect 13556 17580 13562 17644
rect 2606 17440 2922 17441
rect 2606 17376 2612 17440
rect 2676 17376 2692 17440
rect 2756 17376 2772 17440
rect 2836 17376 2852 17440
rect 2916 17376 2922 17440
rect 2606 17375 2922 17376
rect 7606 17440 7922 17441
rect 7606 17376 7612 17440
rect 7676 17376 7692 17440
rect 7756 17376 7772 17440
rect 7836 17376 7852 17440
rect 7916 17376 7922 17440
rect 7606 17375 7922 17376
rect 12606 17440 12922 17441
rect 12606 17376 12612 17440
rect 12676 17376 12692 17440
rect 12756 17376 12772 17440
rect 12836 17376 12852 17440
rect 12916 17376 12922 17440
rect 12606 17375 12922 17376
rect 17606 17440 17922 17441
rect 17606 17376 17612 17440
rect 17676 17376 17692 17440
rect 17756 17376 17772 17440
rect 17836 17376 17852 17440
rect 17916 17376 17922 17440
rect 17606 17375 17922 17376
rect 3877 17370 3943 17373
rect 7465 17370 7531 17373
rect 12433 17370 12499 17373
rect 3877 17368 7531 17370
rect 3877 17312 3882 17368
rect 3938 17312 7470 17368
rect 7526 17312 7531 17368
rect 3877 17310 7531 17312
rect 3877 17307 3943 17310
rect 7465 17307 7531 17310
rect 8894 17368 12499 17370
rect 8894 17312 12438 17368
rect 12494 17312 12499 17368
rect 8894 17310 12499 17312
rect 5349 17234 5415 17237
rect 8894 17234 8954 17310
rect 12433 17307 12499 17310
rect 5349 17232 8954 17234
rect 5349 17176 5354 17232
rect 5410 17176 8954 17232
rect 5349 17174 8954 17176
rect 9121 17234 9187 17237
rect 17309 17234 17375 17237
rect 9121 17232 17375 17234
rect 9121 17176 9126 17232
rect 9182 17176 17314 17232
rect 17370 17176 17375 17232
rect 9121 17174 17375 17176
rect 5349 17171 5415 17174
rect 9121 17171 9187 17174
rect 17309 17171 17375 17174
rect 3366 17036 3372 17100
rect 3436 17098 3442 17100
rect 8661 17098 8727 17101
rect 15142 17098 15148 17100
rect 3436 17038 7436 17098
rect 3436 17036 3442 17038
rect 2405 16964 2471 16965
rect 2405 16960 2452 16964
rect 2516 16962 2522 16964
rect 7376 16962 7436 17038
rect 8661 17096 15148 17098
rect 8661 17040 8666 17096
rect 8722 17040 15148 17096
rect 8661 17038 15148 17040
rect 8661 17035 8727 17038
rect 15142 17036 15148 17038
rect 15212 17036 15218 17100
rect 11513 16962 11579 16965
rect 2405 16904 2410 16960
rect 2405 16900 2452 16904
rect 2516 16902 2562 16962
rect 7376 16960 11579 16962
rect 7376 16904 11518 16960
rect 11574 16904 11579 16960
rect 7376 16902 11579 16904
rect 2516 16900 2522 16902
rect 2405 16899 2471 16900
rect 11513 16899 11579 16902
rect 12341 16962 12407 16965
rect 13905 16962 13971 16965
rect 12341 16960 13971 16962
rect 12341 16904 12346 16960
rect 12402 16904 13910 16960
rect 13966 16904 13971 16960
rect 12341 16902 13971 16904
rect 12341 16899 12407 16902
rect 13905 16899 13971 16902
rect 1946 16896 2262 16897
rect 1946 16832 1952 16896
rect 2016 16832 2032 16896
rect 2096 16832 2112 16896
rect 2176 16832 2192 16896
rect 2256 16832 2262 16896
rect 1946 16831 2262 16832
rect 6946 16896 7262 16897
rect 6946 16832 6952 16896
rect 7016 16832 7032 16896
rect 7096 16832 7112 16896
rect 7176 16832 7192 16896
rect 7256 16832 7262 16896
rect 6946 16831 7262 16832
rect 11946 16896 12262 16897
rect 11946 16832 11952 16896
rect 12016 16832 12032 16896
rect 12096 16832 12112 16896
rect 12176 16832 12192 16896
rect 12256 16832 12262 16896
rect 11946 16831 12262 16832
rect 16946 16896 17262 16897
rect 16946 16832 16952 16896
rect 17016 16832 17032 16896
rect 17096 16832 17112 16896
rect 17176 16832 17192 16896
rect 17256 16832 17262 16896
rect 16946 16831 17262 16832
rect 5441 16828 5507 16829
rect 5390 16826 5396 16828
rect 5350 16766 5396 16826
rect 5460 16824 5507 16828
rect 5502 16768 5507 16824
rect 5390 16764 5396 16766
rect 5460 16764 5507 16768
rect 5441 16763 5507 16764
rect 7465 16826 7531 16829
rect 9070 16826 9076 16828
rect 7465 16824 9076 16826
rect 7465 16768 7470 16824
rect 7526 16768 9076 16824
rect 7465 16766 9076 16768
rect 7465 16763 7531 16766
rect 9070 16764 9076 16766
rect 9140 16764 9146 16828
rect 12433 16826 12499 16829
rect 13302 16826 13308 16828
rect 12433 16824 13308 16826
rect 12433 16768 12438 16824
rect 12494 16768 13308 16824
rect 12433 16766 13308 16768
rect 12433 16763 12499 16766
rect 13302 16764 13308 16766
rect 13372 16764 13378 16828
rect 6310 16628 6316 16692
rect 6380 16690 6386 16692
rect 9121 16690 9187 16693
rect 6380 16688 9187 16690
rect 6380 16632 9126 16688
rect 9182 16632 9187 16688
rect 6380 16630 9187 16632
rect 6380 16628 6386 16630
rect 9121 16627 9187 16630
rect 11329 16690 11395 16693
rect 14549 16690 14615 16693
rect 11329 16688 14615 16690
rect 11329 16632 11334 16688
rect 11390 16632 14554 16688
rect 14610 16632 14615 16688
rect 11329 16630 14615 16632
rect 11329 16627 11395 16630
rect 14549 16627 14615 16630
rect 6545 16554 6611 16557
rect 9857 16554 9923 16557
rect 15193 16554 15259 16557
rect 6545 16552 8218 16554
rect 6545 16496 6550 16552
rect 6606 16496 8218 16552
rect 6545 16494 8218 16496
rect 6545 16491 6611 16494
rect 8158 16418 8218 16494
rect 9857 16552 15259 16554
rect 9857 16496 9862 16552
rect 9918 16496 15198 16552
rect 15254 16496 15259 16552
rect 9857 16494 15259 16496
rect 9857 16491 9923 16494
rect 15193 16491 15259 16494
rect 16614 16492 16620 16556
rect 16684 16554 16690 16556
rect 17125 16554 17191 16557
rect 16684 16552 17191 16554
rect 16684 16496 17130 16552
rect 17186 16496 17191 16552
rect 16684 16494 17191 16496
rect 16684 16492 16690 16494
rect 17125 16491 17191 16494
rect 11789 16418 11855 16421
rect 8158 16416 11855 16418
rect 8158 16360 11794 16416
rect 11850 16360 11855 16416
rect 8158 16358 11855 16360
rect 11789 16355 11855 16358
rect 2606 16352 2922 16353
rect 2606 16288 2612 16352
rect 2676 16288 2692 16352
rect 2756 16288 2772 16352
rect 2836 16288 2852 16352
rect 2916 16288 2922 16352
rect 2606 16287 2922 16288
rect 7606 16352 7922 16353
rect 7606 16288 7612 16352
rect 7676 16288 7692 16352
rect 7756 16288 7772 16352
rect 7836 16288 7852 16352
rect 7916 16288 7922 16352
rect 7606 16287 7922 16288
rect 12606 16352 12922 16353
rect 12606 16288 12612 16352
rect 12676 16288 12692 16352
rect 12756 16288 12772 16352
rect 12836 16288 12852 16352
rect 12916 16288 12922 16352
rect 12606 16287 12922 16288
rect 17606 16352 17922 16353
rect 17606 16288 17612 16352
rect 17676 16288 17692 16352
rect 17756 16288 17772 16352
rect 17836 16288 17852 16352
rect 17916 16288 17922 16352
rect 17606 16287 17922 16288
rect 3693 16282 3759 16285
rect 7465 16282 7531 16285
rect 3693 16280 7531 16282
rect 3693 16224 3698 16280
rect 3754 16224 7470 16280
rect 7526 16224 7531 16280
rect 3693 16222 7531 16224
rect 3693 16219 3759 16222
rect 7465 16219 7531 16222
rect 9438 16220 9444 16284
rect 9508 16282 9514 16284
rect 10593 16282 10659 16285
rect 9508 16280 10659 16282
rect 9508 16224 10598 16280
rect 10654 16224 10659 16280
rect 9508 16222 10659 16224
rect 9508 16220 9514 16222
rect 10593 16219 10659 16222
rect 10726 16220 10732 16284
rect 10796 16282 10802 16284
rect 10796 16222 12450 16282
rect 10796 16220 10802 16222
rect 0 16146 800 16176
rect 1485 16146 1551 16149
rect 0 16144 1551 16146
rect 0 16088 1490 16144
rect 1546 16088 1551 16144
rect 0 16086 1551 16088
rect 0 16056 800 16086
rect 1485 16083 1551 16086
rect 4705 16146 4771 16149
rect 12249 16146 12315 16149
rect 4705 16144 12315 16146
rect 4705 16088 4710 16144
rect 4766 16088 12254 16144
rect 12310 16088 12315 16144
rect 4705 16086 12315 16088
rect 12390 16146 12450 16222
rect 17033 16146 17099 16149
rect 12390 16144 17099 16146
rect 12390 16088 17038 16144
rect 17094 16088 17099 16144
rect 12390 16086 17099 16088
rect 4705 16083 4771 16086
rect 12249 16083 12315 16086
rect 17033 16083 17099 16086
rect 18413 16146 18479 16149
rect 19200 16146 20000 16176
rect 18413 16144 20000 16146
rect 18413 16088 18418 16144
rect 18474 16088 20000 16144
rect 18413 16086 20000 16088
rect 18413 16083 18479 16086
rect 19200 16056 20000 16086
rect 1761 16010 1827 16013
rect 4286 16010 4292 16012
rect 1761 16008 4292 16010
rect 1761 15952 1766 16008
rect 1822 15952 4292 16008
rect 1761 15950 4292 15952
rect 1761 15947 1827 15950
rect 4286 15948 4292 15950
rect 4356 15948 4362 16012
rect 7005 16010 7071 16013
rect 7005 16008 12404 16010
rect 7005 15952 7010 16008
rect 7066 15952 12404 16008
rect 7005 15950 12404 15952
rect 7005 15947 7071 15950
rect 7373 15874 7439 15877
rect 10174 15874 10180 15876
rect 7373 15872 10180 15874
rect 7373 15816 7378 15872
rect 7434 15816 10180 15872
rect 7373 15814 10180 15816
rect 7373 15811 7439 15814
rect 10174 15812 10180 15814
rect 10244 15812 10250 15876
rect 12344 15874 12404 15950
rect 14222 15874 14228 15876
rect 12344 15814 14228 15874
rect 14222 15812 14228 15814
rect 14292 15812 14298 15876
rect 1946 15808 2262 15809
rect 1946 15744 1952 15808
rect 2016 15744 2032 15808
rect 2096 15744 2112 15808
rect 2176 15744 2192 15808
rect 2256 15744 2262 15808
rect 1946 15743 2262 15744
rect 6946 15808 7262 15809
rect 6946 15744 6952 15808
rect 7016 15744 7032 15808
rect 7096 15744 7112 15808
rect 7176 15744 7192 15808
rect 7256 15744 7262 15808
rect 6946 15743 7262 15744
rect 11946 15808 12262 15809
rect 11946 15744 11952 15808
rect 12016 15744 12032 15808
rect 12096 15744 12112 15808
rect 12176 15744 12192 15808
rect 12256 15744 12262 15808
rect 11946 15743 12262 15744
rect 16946 15808 17262 15809
rect 16946 15744 16952 15808
rect 17016 15744 17032 15808
rect 17096 15744 17112 15808
rect 17176 15744 17192 15808
rect 17256 15744 17262 15808
rect 16946 15743 17262 15744
rect 7465 15738 7531 15741
rect 10593 15738 10659 15741
rect 7465 15736 10659 15738
rect 7465 15680 7470 15736
rect 7526 15680 10598 15736
rect 10654 15680 10659 15736
rect 7465 15678 10659 15680
rect 7465 15675 7531 15678
rect 10593 15675 10659 15678
rect 12341 15738 12407 15741
rect 14825 15738 14891 15741
rect 12341 15736 14891 15738
rect 12341 15680 12346 15736
rect 12402 15680 14830 15736
rect 14886 15680 14891 15736
rect 12341 15678 14891 15680
rect 12341 15675 12407 15678
rect 14825 15675 14891 15678
rect 2497 15602 2563 15605
rect 4061 15602 4127 15605
rect 2497 15600 4127 15602
rect 2497 15544 2502 15600
rect 2558 15544 4066 15600
rect 4122 15544 4127 15600
rect 2497 15542 4127 15544
rect 2497 15539 2563 15542
rect 4061 15539 4127 15542
rect 6913 15602 6979 15605
rect 18137 15602 18203 15605
rect 6913 15600 18203 15602
rect 6913 15544 6918 15600
rect 6974 15544 18142 15600
rect 18198 15544 18203 15600
rect 6913 15542 18203 15544
rect 6913 15539 6979 15542
rect 18137 15539 18203 15542
rect 4061 15466 4127 15469
rect 8937 15466 9003 15469
rect 4061 15464 9003 15466
rect 4061 15408 4066 15464
rect 4122 15408 8942 15464
rect 8998 15408 9003 15464
rect 4061 15406 9003 15408
rect 4061 15403 4127 15406
rect 8937 15403 9003 15406
rect 9121 15466 9187 15469
rect 9254 15466 9260 15468
rect 9121 15464 9260 15466
rect 9121 15408 9126 15464
rect 9182 15408 9260 15464
rect 9121 15406 9260 15408
rect 9121 15403 9187 15406
rect 9254 15404 9260 15406
rect 9324 15404 9330 15468
rect 10593 15466 10659 15469
rect 10910 15466 10916 15468
rect 10593 15464 10916 15466
rect 10593 15408 10598 15464
rect 10654 15408 10916 15464
rect 10593 15406 10916 15408
rect 10593 15403 10659 15406
rect 10910 15404 10916 15406
rect 10980 15404 10986 15468
rect 12801 15466 12867 15469
rect 18270 15466 18276 15468
rect 12801 15464 18276 15466
rect 12801 15408 12806 15464
rect 12862 15408 18276 15464
rect 12801 15406 18276 15408
rect 12801 15403 12867 15406
rect 18270 15404 18276 15406
rect 18340 15404 18346 15468
rect 790 15268 796 15332
rect 860 15330 866 15332
rect 1577 15330 1643 15333
rect 860 15328 1643 15330
rect 860 15272 1582 15328
rect 1638 15272 1643 15328
rect 860 15270 1643 15272
rect 860 15268 866 15270
rect 1577 15267 1643 15270
rect 4102 15268 4108 15332
rect 4172 15330 4178 15332
rect 6637 15330 6703 15333
rect 4172 15328 6703 15330
rect 4172 15272 6642 15328
rect 6698 15272 6703 15328
rect 4172 15270 6703 15272
rect 4172 15268 4178 15270
rect 6637 15267 6703 15270
rect 8702 15268 8708 15332
rect 8772 15330 8778 15332
rect 8845 15330 8911 15333
rect 8772 15328 8911 15330
rect 8772 15272 8850 15328
rect 8906 15272 8911 15328
rect 8772 15270 8911 15272
rect 8772 15268 8778 15270
rect 8845 15267 8911 15270
rect 2606 15264 2922 15265
rect 2606 15200 2612 15264
rect 2676 15200 2692 15264
rect 2756 15200 2772 15264
rect 2836 15200 2852 15264
rect 2916 15200 2922 15264
rect 2606 15199 2922 15200
rect 7606 15264 7922 15265
rect 7606 15200 7612 15264
rect 7676 15200 7692 15264
rect 7756 15200 7772 15264
rect 7836 15200 7852 15264
rect 7916 15200 7922 15264
rect 7606 15199 7922 15200
rect 12606 15264 12922 15265
rect 12606 15200 12612 15264
rect 12676 15200 12692 15264
rect 12756 15200 12772 15264
rect 12836 15200 12852 15264
rect 12916 15200 12922 15264
rect 12606 15199 12922 15200
rect 17606 15264 17922 15265
rect 17606 15200 17612 15264
rect 17676 15200 17692 15264
rect 17756 15200 17772 15264
rect 17836 15200 17852 15264
rect 17916 15200 17922 15264
rect 17606 15199 17922 15200
rect 4889 15194 4955 15197
rect 7414 15194 7420 15196
rect 4889 15192 7420 15194
rect 4889 15136 4894 15192
rect 4950 15136 7420 15192
rect 4889 15134 7420 15136
rect 4889 15131 4955 15134
rect 7414 15132 7420 15134
rect 7484 15132 7490 15196
rect 8477 15194 8543 15197
rect 9622 15194 9628 15196
rect 8477 15192 9628 15194
rect 8477 15136 8482 15192
rect 8538 15136 9628 15192
rect 8477 15134 9628 15136
rect 8477 15131 8543 15134
rect 9622 15132 9628 15134
rect 9692 15132 9698 15196
rect 11421 15194 11487 15197
rect 11697 15194 11763 15197
rect 11421 15192 11763 15194
rect 11421 15136 11426 15192
rect 11482 15136 11702 15192
rect 11758 15136 11763 15192
rect 11421 15134 11763 15136
rect 11421 15131 11487 15134
rect 11697 15131 11763 15134
rect 5441 15058 5507 15061
rect 9765 15060 9831 15061
rect 8518 15058 8524 15060
rect 5441 15056 8524 15058
rect 5441 15000 5446 15056
rect 5502 15000 8524 15056
rect 5441 14998 8524 15000
rect 5441 14995 5507 14998
rect 8518 14996 8524 14998
rect 8588 14996 8594 15060
rect 9765 15058 9812 15060
rect 9720 15056 9812 15058
rect 9720 15000 9770 15056
rect 9720 14998 9812 15000
rect 9765 14996 9812 14998
rect 9876 14996 9882 15060
rect 10501 15058 10567 15061
rect 16389 15058 16455 15061
rect 10501 15056 16455 15058
rect 10501 15000 10506 15056
rect 10562 15000 16394 15056
rect 16450 15000 16455 15056
rect 10501 14998 16455 15000
rect 9765 14995 9831 14996
rect 10501 14995 10567 14998
rect 16389 14995 16455 14998
rect 3141 14922 3207 14925
rect 13353 14922 13419 14925
rect 3141 14920 13419 14922
rect 3141 14864 3146 14920
rect 3202 14864 13358 14920
rect 13414 14864 13419 14920
rect 3141 14862 13419 14864
rect 3141 14859 3207 14862
rect 13353 14859 13419 14862
rect 7414 14724 7420 14788
rect 7484 14786 7490 14788
rect 10869 14786 10935 14789
rect 7484 14784 10935 14786
rect 7484 14728 10874 14784
rect 10930 14728 10935 14784
rect 7484 14726 10935 14728
rect 7484 14724 7490 14726
rect 10869 14723 10935 14726
rect 12985 14786 13051 14789
rect 13118 14786 13124 14788
rect 12985 14784 13124 14786
rect 12985 14728 12990 14784
rect 13046 14728 13124 14784
rect 12985 14726 13124 14728
rect 12985 14723 13051 14726
rect 13118 14724 13124 14726
rect 13188 14724 13194 14788
rect 1946 14720 2262 14721
rect 1946 14656 1952 14720
rect 2016 14656 2032 14720
rect 2096 14656 2112 14720
rect 2176 14656 2192 14720
rect 2256 14656 2262 14720
rect 1946 14655 2262 14656
rect 6946 14720 7262 14721
rect 6946 14656 6952 14720
rect 7016 14656 7032 14720
rect 7096 14656 7112 14720
rect 7176 14656 7192 14720
rect 7256 14656 7262 14720
rect 6946 14655 7262 14656
rect 11946 14720 12262 14721
rect 11946 14656 11952 14720
rect 12016 14656 12032 14720
rect 12096 14656 12112 14720
rect 12176 14656 12192 14720
rect 12256 14656 12262 14720
rect 11946 14655 12262 14656
rect 16946 14720 17262 14721
rect 16946 14656 16952 14720
rect 17016 14656 17032 14720
rect 17096 14656 17112 14720
rect 17176 14656 17192 14720
rect 17256 14656 17262 14720
rect 16946 14655 17262 14656
rect 3734 14588 3740 14652
rect 3804 14650 3810 14652
rect 4429 14650 4495 14653
rect 3804 14648 4495 14650
rect 3804 14592 4434 14648
rect 4490 14592 4495 14648
rect 3804 14590 4495 14592
rect 3804 14588 3810 14590
rect 4429 14587 4495 14590
rect 7414 14588 7420 14652
rect 7484 14650 7490 14652
rect 8201 14650 8267 14653
rect 7484 14648 8267 14650
rect 7484 14592 8206 14648
rect 8262 14592 8267 14648
rect 7484 14590 8267 14592
rect 7484 14588 7490 14590
rect 8201 14587 8267 14590
rect 8334 14588 8340 14652
rect 8404 14650 8410 14652
rect 11237 14650 11303 14653
rect 8404 14648 11303 14650
rect 8404 14592 11242 14648
rect 11298 14592 11303 14648
rect 8404 14590 11303 14592
rect 8404 14588 8410 14590
rect 11237 14587 11303 14590
rect 12801 14650 12867 14653
rect 15694 14650 15700 14652
rect 12801 14648 15700 14650
rect 12801 14592 12806 14648
rect 12862 14592 15700 14648
rect 12801 14590 15700 14592
rect 12801 14587 12867 14590
rect 15694 14588 15700 14590
rect 15764 14588 15770 14652
rect 4429 14514 4495 14517
rect 10961 14514 11027 14517
rect 4429 14512 11027 14514
rect 4429 14456 4434 14512
rect 4490 14456 10966 14512
rect 11022 14456 11027 14512
rect 4429 14454 11027 14456
rect 4429 14451 4495 14454
rect 10961 14451 11027 14454
rect 11513 14514 11579 14517
rect 11646 14514 11652 14516
rect 11513 14512 11652 14514
rect 11513 14456 11518 14512
rect 11574 14456 11652 14512
rect 11513 14454 11652 14456
rect 11513 14451 11579 14454
rect 11646 14452 11652 14454
rect 11716 14452 11722 14516
rect 12065 14514 12131 14517
rect 14273 14514 14339 14517
rect 12065 14512 14339 14514
rect 12065 14456 12070 14512
rect 12126 14456 14278 14512
rect 14334 14456 14339 14512
rect 12065 14454 14339 14456
rect 12065 14451 12131 14454
rect 14273 14451 14339 14454
rect 1853 14378 1919 14381
rect 4521 14378 4587 14381
rect 8293 14378 8359 14381
rect 9305 14378 9371 14381
rect 1853 14376 4587 14378
rect 1853 14320 1858 14376
rect 1914 14320 4526 14376
rect 4582 14320 4587 14376
rect 1853 14318 4587 14320
rect 1853 14315 1919 14318
rect 4521 14315 4587 14318
rect 5950 14318 8218 14378
rect 2129 14242 2195 14245
rect 2446 14242 2452 14244
rect 2129 14240 2452 14242
rect 2129 14184 2134 14240
rect 2190 14184 2452 14240
rect 2129 14182 2452 14184
rect 2129 14179 2195 14182
rect 2446 14180 2452 14182
rect 2516 14180 2522 14244
rect 3918 14180 3924 14244
rect 3988 14242 3994 14244
rect 4889 14242 4955 14245
rect 3988 14240 4955 14242
rect 3988 14184 4894 14240
rect 4950 14184 4955 14240
rect 3988 14182 4955 14184
rect 3988 14180 3994 14182
rect 4889 14179 4955 14182
rect 2606 14176 2922 14177
rect 2606 14112 2612 14176
rect 2676 14112 2692 14176
rect 2756 14112 2772 14176
rect 2836 14112 2852 14176
rect 2916 14112 2922 14176
rect 2606 14111 2922 14112
rect 5206 14044 5212 14108
rect 5276 14106 5282 14108
rect 5349 14106 5415 14109
rect 5276 14104 5415 14106
rect 5276 14048 5354 14104
rect 5410 14048 5415 14104
rect 5276 14046 5415 14048
rect 5276 14044 5282 14046
rect 5349 14043 5415 14046
rect 1945 13970 2011 13973
rect 5441 13970 5507 13973
rect 1945 13968 5507 13970
rect 1945 13912 1950 13968
rect 2006 13912 5446 13968
rect 5502 13912 5507 13968
rect 1945 13910 5507 13912
rect 1945 13907 2011 13910
rect 5441 13907 5507 13910
rect 5950 13837 6010 14318
rect 8158 14242 8218 14318
rect 8293 14376 9371 14378
rect 8293 14320 8298 14376
rect 8354 14320 9310 14376
rect 9366 14320 9371 14376
rect 8293 14318 9371 14320
rect 8293 14315 8359 14318
rect 9305 14315 9371 14318
rect 9765 14378 9831 14381
rect 14958 14378 14964 14380
rect 9765 14376 14964 14378
rect 9765 14320 9770 14376
rect 9826 14320 14964 14376
rect 9765 14318 14964 14320
rect 9765 14315 9831 14318
rect 14958 14316 14964 14318
rect 15028 14316 15034 14380
rect 12065 14242 12131 14245
rect 8158 14240 12131 14242
rect 8158 14184 12070 14240
rect 12126 14184 12131 14240
rect 8158 14182 12131 14184
rect 12065 14179 12131 14182
rect 7606 14176 7922 14177
rect 7606 14112 7612 14176
rect 7676 14112 7692 14176
rect 7756 14112 7772 14176
rect 7836 14112 7852 14176
rect 7916 14112 7922 14176
rect 7606 14111 7922 14112
rect 12606 14176 12922 14177
rect 12606 14112 12612 14176
rect 12676 14112 12692 14176
rect 12756 14112 12772 14176
rect 12836 14112 12852 14176
rect 12916 14112 12922 14176
rect 12606 14111 12922 14112
rect 17606 14176 17922 14177
rect 17606 14112 17612 14176
rect 17676 14112 17692 14176
rect 17756 14112 17772 14176
rect 17836 14112 17852 14176
rect 17916 14112 17922 14176
rect 17606 14111 17922 14112
rect 12433 14106 12499 14109
rect 8342 14104 12499 14106
rect 8342 14048 12438 14104
rect 12494 14048 12499 14104
rect 8342 14046 12499 14048
rect 7281 13970 7347 13973
rect 8342 13970 8402 14046
rect 12433 14043 12499 14046
rect 13169 14106 13235 14109
rect 13169 14104 17004 14106
rect 13169 14048 13174 14104
rect 13230 14048 17004 14104
rect 13169 14046 17004 14048
rect 13169 14043 13235 14046
rect 7281 13968 8402 13970
rect 7281 13912 7286 13968
rect 7342 13912 8402 13968
rect 7281 13910 8402 13912
rect 8569 13970 8635 13973
rect 10501 13970 10567 13973
rect 11881 13970 11947 13973
rect 8569 13968 11947 13970
rect 8569 13912 8574 13968
rect 8630 13912 10506 13968
rect 10562 13912 11886 13968
rect 11942 13912 11947 13968
rect 8569 13910 11947 13912
rect 16944 13970 17004 14046
rect 18822 13970 18828 13972
rect 16944 13910 18828 13970
rect 7281 13907 7347 13910
rect 8569 13907 8635 13910
rect 10501 13907 10567 13910
rect 11881 13907 11947 13910
rect 18822 13908 18828 13910
rect 18892 13908 18898 13972
rect 1158 13772 1164 13836
rect 1228 13834 1234 13836
rect 4705 13834 4771 13837
rect 1228 13832 4771 13834
rect 1228 13776 4710 13832
rect 4766 13776 4771 13832
rect 1228 13774 4771 13776
rect 1228 13772 1234 13774
rect 4705 13771 4771 13774
rect 5901 13832 6010 13837
rect 6453 13836 6519 13837
rect 6453 13834 6500 13836
rect 5901 13776 5906 13832
rect 5962 13776 6010 13832
rect 5901 13774 6010 13776
rect 6408 13832 6500 13834
rect 6408 13776 6458 13832
rect 6408 13774 6500 13776
rect 5901 13771 5967 13774
rect 6453 13772 6500 13774
rect 6564 13772 6570 13836
rect 10409 13834 10475 13837
rect 6732 13832 10475 13834
rect 6732 13776 10414 13832
rect 10470 13776 10475 13832
rect 6732 13774 10475 13776
rect 6453 13771 6519 13772
rect 0 13698 800 13728
rect 1485 13698 1551 13701
rect 0 13696 1551 13698
rect 0 13640 1490 13696
rect 1546 13640 1551 13696
rect 0 13638 1551 13640
rect 0 13608 800 13638
rect 1485 13635 1551 13638
rect 3182 13636 3188 13700
rect 3252 13698 3258 13700
rect 6732 13698 6792 13774
rect 10409 13771 10475 13774
rect 11421 13834 11487 13837
rect 13445 13834 13511 13837
rect 11421 13832 13511 13834
rect 11421 13776 11426 13832
rect 11482 13776 13450 13832
rect 13506 13776 13511 13832
rect 11421 13774 13511 13776
rect 11421 13771 11487 13774
rect 13445 13771 13511 13774
rect 14733 13834 14799 13837
rect 16614 13834 16620 13836
rect 14733 13832 16620 13834
rect 14733 13776 14738 13832
rect 14794 13776 16620 13832
rect 14733 13774 16620 13776
rect 14733 13771 14799 13774
rect 16614 13772 16620 13774
rect 16684 13772 16690 13836
rect 3252 13638 6792 13698
rect 3252 13636 3258 13638
rect 8518 13636 8524 13700
rect 8588 13698 8594 13700
rect 11462 13698 11468 13700
rect 8588 13638 11468 13698
rect 8588 13636 8594 13638
rect 11462 13636 11468 13638
rect 11532 13636 11538 13700
rect 18413 13698 18479 13701
rect 19200 13698 20000 13728
rect 18413 13696 20000 13698
rect 18413 13640 18418 13696
rect 18474 13640 20000 13696
rect 18413 13638 20000 13640
rect 18413 13635 18479 13638
rect 1946 13632 2262 13633
rect 1946 13568 1952 13632
rect 2016 13568 2032 13632
rect 2096 13568 2112 13632
rect 2176 13568 2192 13632
rect 2256 13568 2262 13632
rect 1946 13567 2262 13568
rect 6946 13632 7262 13633
rect 6946 13568 6952 13632
rect 7016 13568 7032 13632
rect 7096 13568 7112 13632
rect 7176 13568 7192 13632
rect 7256 13568 7262 13632
rect 6946 13567 7262 13568
rect 11946 13632 12262 13633
rect 11946 13568 11952 13632
rect 12016 13568 12032 13632
rect 12096 13568 12112 13632
rect 12176 13568 12192 13632
rect 12256 13568 12262 13632
rect 11946 13567 12262 13568
rect 16946 13632 17262 13633
rect 16946 13568 16952 13632
rect 17016 13568 17032 13632
rect 17096 13568 17112 13632
rect 17176 13568 17192 13632
rect 17256 13568 17262 13632
rect 19200 13608 20000 13638
rect 16946 13567 17262 13568
rect 4061 13562 4127 13565
rect 5533 13562 5599 13565
rect 5758 13562 5764 13564
rect 2454 13560 4127 13562
rect 2454 13504 4066 13560
rect 4122 13504 4127 13560
rect 2454 13502 4127 13504
rect 1342 13364 1348 13428
rect 1412 13426 1418 13428
rect 2454 13426 2514 13502
rect 4061 13499 4127 13502
rect 4294 13560 5764 13562
rect 4294 13504 5538 13560
rect 5594 13504 5764 13560
rect 4294 13502 5764 13504
rect 1412 13366 2514 13426
rect 1412 13364 1418 13366
rect 2998 13364 3004 13428
rect 3068 13426 3074 13428
rect 4294 13426 4354 13502
rect 5533 13499 5599 13502
rect 5758 13500 5764 13502
rect 5828 13500 5834 13564
rect 5942 13500 5948 13564
rect 6012 13562 6018 13564
rect 6085 13562 6151 13565
rect 6012 13560 6151 13562
rect 6012 13504 6090 13560
rect 6146 13504 6151 13560
rect 6012 13502 6151 13504
rect 6012 13500 6018 13502
rect 6085 13499 6151 13502
rect 6453 13562 6519 13565
rect 6678 13562 6684 13564
rect 6453 13560 6684 13562
rect 6453 13504 6458 13560
rect 6514 13504 6684 13560
rect 6453 13502 6684 13504
rect 6453 13499 6519 13502
rect 6678 13500 6684 13502
rect 6748 13500 6754 13564
rect 7925 13562 7991 13565
rect 11697 13562 11763 13565
rect 7925 13560 11763 13562
rect 7925 13504 7930 13560
rect 7986 13504 11702 13560
rect 11758 13504 11763 13560
rect 7925 13502 11763 13504
rect 7925 13499 7991 13502
rect 11697 13499 11763 13502
rect 17493 13562 17559 13565
rect 18638 13562 18644 13564
rect 17493 13560 18644 13562
rect 17493 13504 17498 13560
rect 17554 13504 18644 13560
rect 17493 13502 18644 13504
rect 17493 13499 17559 13502
rect 18638 13500 18644 13502
rect 18708 13500 18714 13564
rect 3068 13366 4354 13426
rect 3068 13364 3074 13366
rect 4838 13364 4844 13428
rect 4908 13426 4914 13428
rect 4981 13426 5047 13429
rect 8293 13426 8359 13429
rect 4908 13424 8359 13426
rect 4908 13368 4986 13424
rect 5042 13368 8298 13424
rect 8354 13368 8359 13424
rect 4908 13366 8359 13368
rect 4908 13364 4914 13366
rect 4981 13363 5047 13366
rect 8293 13363 8359 13366
rect 9990 13364 9996 13428
rect 10060 13426 10066 13428
rect 10133 13426 10199 13429
rect 10060 13424 10199 13426
rect 10060 13368 10138 13424
rect 10194 13368 10199 13424
rect 10060 13366 10199 13368
rect 10060 13364 10066 13366
rect 10133 13363 10199 13366
rect 10542 13364 10548 13428
rect 10612 13426 10618 13428
rect 14181 13426 14247 13429
rect 10612 13424 14247 13426
rect 10612 13368 14186 13424
rect 14242 13368 14247 13424
rect 10612 13366 14247 13368
rect 10612 13364 10618 13366
rect 14181 13363 14247 13366
rect 2865 13290 2931 13293
rect 5809 13290 5875 13293
rect 2865 13288 5875 13290
rect 2865 13232 2870 13288
rect 2926 13232 5814 13288
rect 5870 13232 5875 13288
rect 2865 13230 5875 13232
rect 2865 13227 2931 13230
rect 5809 13227 5875 13230
rect 6177 13290 6243 13293
rect 7189 13290 7255 13293
rect 7557 13290 7623 13293
rect 6177 13288 7255 13290
rect 6177 13232 6182 13288
rect 6238 13232 7194 13288
rect 7250 13232 7255 13288
rect 6177 13230 7255 13232
rect 6177 13227 6243 13230
rect 7189 13227 7255 13230
rect 7376 13288 7623 13290
rect 7376 13232 7562 13288
rect 7618 13232 7623 13288
rect 7376 13230 7623 13232
rect 7376 13157 7436 13230
rect 7557 13227 7623 13230
rect 7741 13290 7807 13293
rect 8569 13290 8635 13293
rect 7741 13288 8635 13290
rect 7741 13232 7746 13288
rect 7802 13232 8574 13288
rect 8630 13232 8635 13288
rect 7741 13230 8635 13232
rect 7741 13227 7807 13230
rect 8569 13227 8635 13230
rect 9213 13290 9279 13293
rect 10358 13290 10364 13292
rect 9213 13288 10364 13290
rect 9213 13232 9218 13288
rect 9274 13232 10364 13288
rect 9213 13230 10364 13232
rect 9213 13227 9279 13230
rect 10358 13228 10364 13230
rect 10428 13228 10434 13292
rect 11094 13228 11100 13292
rect 11164 13290 11170 13292
rect 11237 13290 11303 13293
rect 15469 13290 15535 13293
rect 11164 13288 11303 13290
rect 11164 13232 11242 13288
rect 11298 13232 11303 13288
rect 11164 13230 11303 13232
rect 11164 13228 11170 13230
rect 11237 13227 11303 13230
rect 11424 13288 15535 13290
rect 11424 13232 15474 13288
rect 15530 13232 15535 13288
rect 11424 13230 15535 13232
rect 4245 13154 4311 13157
rect 7373 13154 7439 13157
rect 4245 13152 7439 13154
rect 4245 13096 4250 13152
rect 4306 13096 7378 13152
rect 7434 13096 7439 13152
rect 4245 13094 7439 13096
rect 4245 13091 4311 13094
rect 7373 13091 7439 13094
rect 8477 13156 8543 13157
rect 8477 13152 8524 13156
rect 8588 13154 8594 13156
rect 8477 13096 8482 13152
rect 8477 13092 8524 13096
rect 8588 13094 8634 13154
rect 8588 13092 8594 13094
rect 9070 13092 9076 13156
rect 9140 13154 9146 13156
rect 9305 13154 9371 13157
rect 9806 13154 9812 13156
rect 9140 13152 9371 13154
rect 9140 13096 9310 13152
rect 9366 13096 9371 13152
rect 9140 13094 9371 13096
rect 9140 13092 9146 13094
rect 8477 13091 8543 13092
rect 9305 13091 9371 13094
rect 9446 13094 9812 13154
rect 2606 13088 2922 13089
rect 2606 13024 2612 13088
rect 2676 13024 2692 13088
rect 2756 13024 2772 13088
rect 2836 13024 2852 13088
rect 2916 13024 2922 13088
rect 2606 13023 2922 13024
rect 7606 13088 7922 13089
rect 7606 13024 7612 13088
rect 7676 13024 7692 13088
rect 7756 13024 7772 13088
rect 7836 13024 7852 13088
rect 7916 13024 7922 13088
rect 7606 13023 7922 13024
rect 3233 13018 3299 13021
rect 3233 13016 3618 13018
rect 3233 12960 3238 13016
rect 3294 12960 3618 13016
rect 3233 12958 3618 12960
rect 3233 12955 3299 12958
rect 2957 12882 3023 12885
rect 3325 12882 3391 12885
rect 2957 12880 3391 12882
rect 2957 12824 2962 12880
rect 3018 12824 3330 12880
rect 3386 12824 3391 12880
rect 2957 12822 3391 12824
rect 3558 12882 3618 12958
rect 4654 12956 4660 13020
rect 4724 13018 4730 13020
rect 5625 13018 5691 13021
rect 4724 13016 5691 13018
rect 4724 12960 5630 13016
rect 5686 12960 5691 13016
rect 4724 12958 5691 12960
rect 4724 12956 4730 12958
rect 5625 12955 5691 12958
rect 6361 13018 6427 13021
rect 7281 13018 7347 13021
rect 6361 13016 7347 13018
rect 6361 12960 6366 13016
rect 6422 12960 7286 13016
rect 7342 12960 7347 13016
rect 6361 12958 7347 12960
rect 6361 12955 6427 12958
rect 7281 12955 7347 12958
rect 9070 12956 9076 13020
rect 9140 13018 9146 13020
rect 9446 13018 9506 13094
rect 9806 13092 9812 13094
rect 9876 13154 9882 13156
rect 11424 13154 11484 13230
rect 15469 13227 15535 13230
rect 9876 13094 11484 13154
rect 9876 13092 9882 13094
rect 12606 13088 12922 13089
rect 12606 13024 12612 13088
rect 12676 13024 12692 13088
rect 12756 13024 12772 13088
rect 12836 13024 12852 13088
rect 12916 13024 12922 13088
rect 12606 13023 12922 13024
rect 17606 13088 17922 13089
rect 17606 13024 17612 13088
rect 17676 13024 17692 13088
rect 17756 13024 17772 13088
rect 17836 13024 17852 13088
rect 17916 13024 17922 13088
rect 17606 13023 17922 13024
rect 9140 12958 9506 13018
rect 9857 13018 9923 13021
rect 10542 13018 10548 13020
rect 9857 13016 10548 13018
rect 9857 12960 9862 13016
rect 9918 12960 10548 13016
rect 9857 12958 10548 12960
rect 9140 12956 9146 12958
rect 9857 12955 9923 12958
rect 10542 12956 10548 12958
rect 10612 12956 10618 13020
rect 10777 13018 10843 13021
rect 11237 13018 11303 13021
rect 10777 13016 11303 13018
rect 10777 12960 10782 13016
rect 10838 12960 11242 13016
rect 11298 12960 11303 13016
rect 10777 12958 11303 12960
rect 10777 12955 10843 12958
rect 11237 12955 11303 12958
rect 13077 13018 13143 13021
rect 16297 13018 16363 13021
rect 13077 13016 16363 13018
rect 13077 12960 13082 13016
rect 13138 12960 16302 13016
rect 16358 12960 16363 13016
rect 13077 12958 16363 12960
rect 13077 12955 13143 12958
rect 16297 12955 16363 12958
rect 6177 12882 6243 12885
rect 3558 12880 6243 12882
rect 3558 12824 6182 12880
rect 6238 12824 6243 12880
rect 3558 12822 6243 12824
rect 2957 12819 3023 12822
rect 3325 12819 3391 12822
rect 6177 12819 6243 12822
rect 6545 12882 6611 12885
rect 9673 12882 9739 12885
rect 6545 12880 9739 12882
rect 6545 12824 6550 12880
rect 6606 12824 9678 12880
rect 9734 12824 9739 12880
rect 6545 12822 9739 12824
rect 6545 12819 6611 12822
rect 9673 12819 9739 12822
rect 10133 12882 10199 12885
rect 10593 12882 10659 12885
rect 10133 12880 10659 12882
rect 10133 12824 10138 12880
rect 10194 12824 10598 12880
rect 10654 12824 10659 12880
rect 10133 12822 10659 12824
rect 10133 12819 10199 12822
rect 10593 12819 10659 12822
rect 10869 12882 10935 12885
rect 11053 12882 11119 12885
rect 10869 12880 11119 12882
rect 10869 12824 10874 12880
rect 10930 12824 11058 12880
rect 11114 12824 11119 12880
rect 10869 12822 11119 12824
rect 10869 12819 10935 12822
rect 11053 12819 11119 12822
rect 11697 12882 11763 12885
rect 17677 12882 17743 12885
rect 11697 12880 17743 12882
rect 11697 12824 11702 12880
rect 11758 12824 17682 12880
rect 17738 12824 17743 12880
rect 11697 12822 17743 12824
rect 11697 12819 11763 12822
rect 17677 12819 17743 12822
rect 18229 12882 18295 12885
rect 19006 12882 19012 12884
rect 18229 12880 19012 12882
rect 18229 12824 18234 12880
rect 18290 12824 19012 12880
rect 18229 12822 19012 12824
rect 18229 12819 18295 12822
rect 19006 12820 19012 12822
rect 19076 12820 19082 12884
rect 2773 12746 2839 12749
rect 6545 12746 6611 12749
rect 2773 12744 6611 12746
rect 2773 12688 2778 12744
rect 2834 12688 6550 12744
rect 6606 12688 6611 12744
rect 2773 12686 6611 12688
rect 2773 12683 2839 12686
rect 6545 12683 6611 12686
rect 6729 12746 6795 12749
rect 9765 12748 9831 12749
rect 8886 12746 8892 12748
rect 6729 12744 8892 12746
rect 6729 12688 6734 12744
rect 6790 12688 8892 12744
rect 6729 12686 8892 12688
rect 6729 12683 6795 12686
rect 8886 12684 8892 12686
rect 8956 12684 8962 12748
rect 9765 12744 9812 12748
rect 9876 12746 9882 12748
rect 11329 12746 11395 12749
rect 9765 12688 9770 12744
rect 9765 12684 9812 12688
rect 9876 12686 10242 12746
rect 9876 12684 9882 12686
rect 9765 12683 9831 12684
rect 2865 12610 2931 12613
rect 4337 12610 4403 12613
rect 6361 12610 6427 12613
rect 2865 12608 6427 12610
rect 2865 12552 2870 12608
rect 2926 12552 4342 12608
rect 4398 12552 6366 12608
rect 6422 12552 6427 12608
rect 2865 12550 6427 12552
rect 2865 12547 2931 12550
rect 4337 12547 4403 12550
rect 6361 12547 6427 12550
rect 7465 12610 7531 12613
rect 9949 12610 10015 12613
rect 7465 12608 10015 12610
rect 7465 12552 7470 12608
rect 7526 12552 9954 12608
rect 10010 12552 10015 12608
rect 7465 12550 10015 12552
rect 10182 12610 10242 12686
rect 10550 12744 11395 12746
rect 10550 12688 11334 12744
rect 11390 12688 11395 12744
rect 10550 12686 11395 12688
rect 10550 12610 10610 12686
rect 11329 12683 11395 12686
rect 11605 12746 11671 12749
rect 17677 12746 17743 12749
rect 11605 12744 17743 12746
rect 11605 12688 11610 12744
rect 11666 12688 17682 12744
rect 17738 12688 17743 12744
rect 11605 12686 17743 12688
rect 11605 12683 11671 12686
rect 17677 12683 17743 12686
rect 10182 12550 10610 12610
rect 7465 12547 7531 12550
rect 9949 12547 10015 12550
rect 10910 12548 10916 12612
rect 10980 12610 10986 12612
rect 11513 12610 11579 12613
rect 10980 12608 11579 12610
rect 10980 12552 11518 12608
rect 11574 12552 11579 12608
rect 10980 12550 11579 12552
rect 10980 12548 10986 12550
rect 11513 12547 11579 12550
rect 15653 12610 15719 12613
rect 15929 12610 15995 12613
rect 15653 12608 15995 12610
rect 15653 12552 15658 12608
rect 15714 12552 15934 12608
rect 15990 12552 15995 12608
rect 15653 12550 15995 12552
rect 15653 12547 15719 12550
rect 15929 12547 15995 12550
rect 1946 12544 2262 12545
rect 1946 12480 1952 12544
rect 2016 12480 2032 12544
rect 2096 12480 2112 12544
rect 2176 12480 2192 12544
rect 2256 12480 2262 12544
rect 1946 12479 2262 12480
rect 6946 12544 7262 12545
rect 6946 12480 6952 12544
rect 7016 12480 7032 12544
rect 7096 12480 7112 12544
rect 7176 12480 7192 12544
rect 7256 12480 7262 12544
rect 6946 12479 7262 12480
rect 11946 12544 12262 12545
rect 11946 12480 11952 12544
rect 12016 12480 12032 12544
rect 12096 12480 12112 12544
rect 12176 12480 12192 12544
rect 12256 12480 12262 12544
rect 11946 12479 12262 12480
rect 16946 12544 17262 12545
rect 16946 12480 16952 12544
rect 17016 12480 17032 12544
rect 17096 12480 17112 12544
rect 17176 12480 17192 12544
rect 17256 12480 17262 12544
rect 16946 12479 17262 12480
rect 3417 12474 3483 12477
rect 3877 12474 3943 12477
rect 4613 12474 4679 12477
rect 10593 12474 10659 12477
rect 11789 12474 11855 12477
rect 3417 12472 3943 12474
rect 1025 12450 1091 12453
rect 982 12448 1091 12450
rect 982 12392 1030 12448
rect 1086 12392 1091 12448
rect 3417 12416 3422 12472
rect 3478 12416 3882 12472
rect 3938 12416 3943 12472
rect 3417 12414 3943 12416
rect 3417 12411 3483 12414
rect 3877 12411 3943 12414
rect 4110 12472 6746 12474
rect 4110 12416 4618 12472
rect 4674 12416 6746 12472
rect 4110 12414 6746 12416
rect 982 12387 1091 12392
rect 105 12338 171 12341
rect 982 12338 1042 12387
rect 4110 12338 4170 12414
rect 4613 12411 4679 12414
rect 105 12336 1042 12338
rect 105 12280 110 12336
rect 166 12280 1042 12336
rect 105 12278 1042 12280
rect 1350 12278 4170 12338
rect 4613 12338 4679 12341
rect 5809 12340 5875 12341
rect 5022 12338 5028 12340
rect 4613 12336 5028 12338
rect 4613 12280 4618 12336
rect 4674 12280 5028 12336
rect 4613 12278 5028 12280
rect 105 12275 171 12278
rect 1209 12202 1275 12205
rect 1350 12202 1410 12278
rect 4613 12275 4679 12278
rect 5022 12276 5028 12278
rect 5092 12276 5098 12340
rect 5758 12338 5764 12340
rect 5718 12278 5764 12338
rect 5828 12336 5875 12340
rect 5870 12280 5875 12336
rect 5758 12276 5764 12278
rect 5828 12276 5875 12280
rect 6686 12338 6746 12414
rect 7422 12472 10659 12474
rect 7422 12416 10598 12472
rect 10654 12416 10659 12472
rect 7422 12414 10659 12416
rect 7422 12338 7482 12414
rect 10593 12411 10659 12414
rect 10734 12472 11855 12474
rect 10734 12416 11794 12472
rect 11850 12416 11855 12472
rect 10734 12414 11855 12416
rect 6686 12278 7482 12338
rect 7649 12338 7715 12341
rect 10734 12338 10794 12414
rect 11789 12411 11855 12414
rect 14273 12338 14339 12341
rect 14549 12338 14615 12341
rect 7649 12336 10794 12338
rect 7649 12280 7654 12336
rect 7710 12280 10794 12336
rect 7649 12278 10794 12280
rect 10872 12278 13508 12338
rect 5809 12275 5875 12276
rect 7649 12275 7715 12278
rect 1209 12200 1410 12202
rect 1209 12144 1214 12200
rect 1270 12144 1410 12200
rect 1209 12142 1410 12144
rect 2589 12202 2655 12205
rect 6361 12202 6427 12205
rect 7097 12202 7163 12205
rect 9949 12202 10015 12205
rect 2589 12200 7163 12202
rect 2589 12144 2594 12200
rect 2650 12144 6366 12200
rect 6422 12144 7102 12200
rect 7158 12144 7163 12200
rect 2589 12142 7163 12144
rect 1209 12139 1275 12142
rect 2589 12139 2655 12142
rect 6361 12139 6427 12142
rect 7097 12139 7163 12142
rect 7238 12200 10015 12202
rect 7238 12144 9954 12200
rect 10010 12144 10015 12200
rect 7238 12142 10015 12144
rect 3785 12066 3851 12069
rect 7238 12066 7298 12142
rect 9949 12139 10015 12142
rect 3785 12064 7298 12066
rect 3785 12008 3790 12064
rect 3846 12008 7298 12064
rect 3785 12006 7298 12008
rect 3785 12003 3851 12006
rect 8150 12004 8156 12068
rect 8220 12066 8226 12068
rect 9254 12066 9260 12068
rect 8220 12006 9260 12066
rect 8220 12004 8226 12006
rect 9254 12004 9260 12006
rect 9324 12004 9330 12068
rect 9673 12066 9739 12069
rect 10872 12066 10932 12278
rect 11278 12140 11284 12204
rect 11348 12202 11354 12204
rect 12382 12202 12388 12204
rect 11348 12142 12388 12202
rect 11348 12140 11354 12142
rect 12382 12140 12388 12142
rect 12452 12140 12458 12204
rect 12985 12200 13051 12205
rect 12985 12144 12990 12200
rect 13046 12144 13051 12200
rect 12985 12139 13051 12144
rect 13169 12202 13235 12205
rect 13302 12202 13308 12204
rect 13169 12200 13308 12202
rect 13169 12144 13174 12200
rect 13230 12144 13308 12200
rect 13169 12142 13308 12144
rect 13169 12139 13235 12142
rect 13302 12140 13308 12142
rect 13372 12140 13378 12204
rect 9673 12064 10932 12066
rect 9673 12008 9678 12064
rect 9734 12008 10932 12064
rect 9673 12006 10932 12008
rect 9673 12003 9739 12006
rect 2606 12000 2922 12001
rect 2606 11936 2612 12000
rect 2676 11936 2692 12000
rect 2756 11936 2772 12000
rect 2836 11936 2852 12000
rect 2916 11936 2922 12000
rect 2606 11935 2922 11936
rect 7606 12000 7922 12001
rect 7606 11936 7612 12000
rect 7676 11936 7692 12000
rect 7756 11936 7772 12000
rect 7836 11936 7852 12000
rect 7916 11936 7922 12000
rect 7606 11935 7922 11936
rect 12606 12000 12922 12001
rect 12606 11936 12612 12000
rect 12676 11936 12692 12000
rect 12756 11936 12772 12000
rect 12836 11936 12852 12000
rect 12916 11936 12922 12000
rect 12606 11935 12922 11936
rect 3601 11930 3667 11933
rect 8017 11930 8083 11933
rect 12433 11930 12499 11933
rect 3601 11928 6792 11930
rect 3601 11872 3606 11928
rect 3662 11872 6792 11928
rect 3601 11870 6792 11872
rect 3601 11867 3667 11870
rect 4061 11794 4127 11797
rect 4245 11794 4311 11797
rect 4061 11792 4311 11794
rect 4061 11736 4066 11792
rect 4122 11736 4250 11792
rect 4306 11736 4311 11792
rect 4061 11734 4311 11736
rect 4061 11731 4127 11734
rect 4245 11731 4311 11734
rect 4797 11794 4863 11797
rect 5022 11794 5028 11796
rect 4797 11792 5028 11794
rect 4797 11736 4802 11792
rect 4858 11736 5028 11792
rect 4797 11734 5028 11736
rect 4797 11731 4863 11734
rect 5022 11732 5028 11734
rect 5092 11732 5098 11796
rect 5349 11794 5415 11797
rect 5993 11794 6059 11797
rect 5349 11792 6059 11794
rect 5349 11736 5354 11792
rect 5410 11736 5998 11792
rect 6054 11736 6059 11792
rect 5349 11734 6059 11736
rect 5349 11731 5415 11734
rect 5993 11731 6059 11734
rect 6732 11794 6792 11870
rect 8017 11928 12499 11930
rect 8017 11872 8022 11928
rect 8078 11872 12438 11928
rect 12494 11872 12499 11928
rect 8017 11870 12499 11872
rect 12988 11930 13048 12139
rect 13448 12066 13508 12278
rect 14273 12336 14615 12338
rect 14273 12280 14278 12336
rect 14334 12280 14554 12336
rect 14610 12280 14615 12336
rect 14273 12278 14615 12280
rect 14273 12275 14339 12278
rect 14549 12275 14615 12278
rect 15142 12276 15148 12340
rect 15212 12338 15218 12340
rect 15212 12278 16682 12338
rect 15212 12276 15218 12278
rect 13670 12140 13676 12204
rect 13740 12202 13746 12204
rect 14181 12202 14247 12205
rect 13740 12200 14247 12202
rect 13740 12144 14186 12200
rect 14242 12144 14247 12200
rect 13740 12142 14247 12144
rect 13740 12140 13746 12142
rect 14181 12139 14247 12142
rect 15142 12140 15148 12204
rect 15212 12202 15218 12204
rect 16481 12202 16547 12205
rect 15212 12200 16547 12202
rect 15212 12144 16486 12200
rect 16542 12144 16547 12200
rect 15212 12142 16547 12144
rect 16622 12202 16682 12278
rect 18454 12202 18460 12204
rect 16622 12142 18460 12202
rect 15212 12140 15218 12142
rect 16481 12139 16547 12142
rect 18454 12140 18460 12142
rect 18524 12140 18530 12204
rect 14273 12066 14339 12069
rect 13448 12064 14339 12066
rect 13448 12008 14278 12064
rect 14334 12008 14339 12064
rect 13448 12006 14339 12008
rect 14273 12003 14339 12006
rect 17606 12000 17922 12001
rect 17606 11936 17612 12000
rect 17676 11936 17692 12000
rect 17756 11936 17772 12000
rect 17836 11936 17852 12000
rect 17916 11936 17922 12000
rect 17606 11935 17922 11936
rect 13997 11930 14063 11933
rect 12988 11928 14063 11930
rect 12988 11872 14002 11928
rect 14058 11872 14063 11928
rect 12988 11870 14063 11872
rect 8017 11867 8083 11870
rect 12433 11867 12499 11870
rect 13997 11867 14063 11870
rect 16246 11868 16252 11932
rect 16316 11930 16322 11932
rect 17401 11930 17467 11933
rect 16316 11928 17467 11930
rect 16316 11872 17406 11928
rect 17462 11872 17467 11928
rect 16316 11870 17467 11872
rect 16316 11868 16322 11870
rect 17401 11867 17467 11870
rect 10869 11796 10935 11797
rect 6732 11734 10012 11794
rect 1485 11658 1551 11661
rect 5901 11658 5967 11661
rect 1485 11656 5967 11658
rect 1485 11600 1490 11656
rect 1546 11600 5906 11656
rect 5962 11600 5967 11656
rect 1485 11598 5967 11600
rect 1485 11595 1551 11598
rect 5901 11595 5967 11598
rect 6732 11525 6792 11734
rect 7097 11658 7163 11661
rect 9765 11658 9831 11661
rect 7097 11656 9831 11658
rect 7097 11600 7102 11656
rect 7158 11600 9770 11656
rect 9826 11600 9831 11656
rect 7097 11598 9831 11600
rect 9952 11658 10012 11734
rect 10174 11732 10180 11796
rect 10244 11794 10250 11796
rect 10869 11794 10916 11796
rect 10244 11792 10916 11794
rect 10244 11736 10874 11792
rect 10244 11734 10916 11736
rect 10244 11732 10250 11734
rect 10869 11732 10916 11734
rect 10980 11732 10986 11796
rect 11789 11794 11855 11797
rect 16665 11794 16731 11797
rect 11789 11792 16731 11794
rect 11789 11736 11794 11792
rect 11850 11736 16670 11792
rect 16726 11736 16731 11792
rect 11789 11734 16731 11736
rect 10869 11731 10935 11732
rect 11789 11731 11855 11734
rect 16665 11731 16731 11734
rect 18321 11658 18387 11661
rect 9952 11656 18387 11658
rect 9952 11600 18326 11656
rect 18382 11600 18387 11656
rect 9952 11598 18387 11600
rect 7097 11595 7163 11598
rect 9765 11595 9831 11598
rect 18321 11595 18387 11598
rect 2446 11460 2452 11524
rect 2516 11522 2522 11524
rect 6177 11522 6243 11525
rect 2516 11520 6243 11522
rect 2516 11464 6182 11520
rect 6238 11464 6243 11520
rect 2516 11462 6243 11464
rect 2516 11460 2522 11462
rect 6177 11459 6243 11462
rect 6729 11520 6795 11525
rect 6729 11464 6734 11520
rect 6790 11464 6795 11520
rect 6729 11459 6795 11464
rect 7373 11522 7439 11525
rect 9673 11522 9739 11525
rect 7373 11520 9739 11522
rect 7373 11464 7378 11520
rect 7434 11464 9678 11520
rect 9734 11464 9739 11520
rect 7373 11462 9739 11464
rect 7373 11459 7439 11462
rect 9673 11459 9739 11462
rect 9949 11522 10015 11525
rect 13261 11522 13327 11525
rect 13905 11522 13971 11525
rect 9949 11520 11162 11522
rect 9949 11464 9954 11520
rect 10010 11464 11162 11520
rect 9949 11462 11162 11464
rect 9949 11459 10015 11462
rect 1946 11456 2262 11457
rect 1946 11392 1952 11456
rect 2016 11392 2032 11456
rect 2096 11392 2112 11456
rect 2176 11392 2192 11456
rect 2256 11392 2262 11456
rect 1946 11391 2262 11392
rect 6946 11456 7262 11457
rect 6946 11392 6952 11456
rect 7016 11392 7032 11456
rect 7096 11392 7112 11456
rect 7176 11392 7192 11456
rect 7256 11392 7262 11456
rect 6946 11391 7262 11392
rect 4429 11388 4495 11389
rect 4429 11384 4476 11388
rect 4540 11386 4546 11388
rect 4705 11386 4771 11389
rect 5073 11386 5139 11389
rect 5717 11386 5783 11389
rect 4429 11328 4434 11384
rect 4429 11324 4476 11328
rect 4540 11326 4586 11386
rect 4705 11384 5783 11386
rect 4705 11328 4710 11384
rect 4766 11328 5078 11384
rect 5134 11328 5722 11384
rect 5778 11328 5783 11384
rect 4705 11326 5783 11328
rect 4540 11324 4546 11326
rect 4429 11323 4495 11324
rect 4705 11323 4771 11326
rect 5073 11323 5139 11326
rect 5717 11323 5783 11326
rect 7925 11386 7991 11389
rect 9213 11388 9279 11389
rect 8334 11386 8340 11388
rect 7925 11384 8340 11386
rect 7925 11328 7930 11384
rect 7986 11328 8340 11384
rect 7925 11326 8340 11328
rect 7925 11323 7991 11326
rect 8334 11324 8340 11326
rect 8404 11324 8410 11388
rect 9213 11386 9260 11388
rect 9168 11384 9260 11386
rect 9168 11328 9218 11384
rect 9168 11326 9260 11328
rect 9213 11324 9260 11326
rect 9324 11324 9330 11388
rect 9622 11324 9628 11388
rect 9692 11386 9698 11388
rect 10961 11386 11027 11389
rect 9692 11384 11027 11386
rect 9692 11328 10966 11384
rect 11022 11328 11027 11384
rect 9692 11326 11027 11328
rect 9692 11324 9698 11326
rect 9213 11323 9279 11324
rect 10961 11323 11027 11326
rect 0 11250 800 11280
rect 1393 11250 1459 11253
rect 4613 11252 4679 11253
rect 4613 11250 4660 11252
rect 0 11248 1459 11250
rect 0 11192 1398 11248
rect 1454 11192 1459 11248
rect 0 11190 1459 11192
rect 4568 11248 4660 11250
rect 4568 11192 4618 11248
rect 4568 11190 4660 11192
rect 0 11160 800 11190
rect 1393 11187 1459 11190
rect 4613 11188 4660 11190
rect 4724 11188 4730 11252
rect 5574 11188 5580 11252
rect 5644 11250 5650 11252
rect 5809 11250 5875 11253
rect 5644 11248 5875 11250
rect 5644 11192 5814 11248
rect 5870 11192 5875 11248
rect 5644 11190 5875 11192
rect 5644 11188 5650 11190
rect 4613 11187 4679 11188
rect 5809 11187 5875 11190
rect 6824 11250 7344 11284
rect 7925 11250 7991 11253
rect 9216 11250 9276 11323
rect 10964 11253 11024 11323
rect 6824 11224 7436 11250
rect 5073 11114 5139 11117
rect 6824 11114 6884 11224
rect 7284 11190 7436 11224
rect 2454 11054 3066 11114
rect 1117 10978 1183 10981
rect 2454 10978 2514 11054
rect 1117 10976 2514 10978
rect 1117 10920 1122 10976
rect 1178 10920 2514 10976
rect 1117 10918 2514 10920
rect 3006 10978 3066 11054
rect 5073 11112 6884 11114
rect 5073 11056 5078 11112
rect 5134 11056 6884 11112
rect 5073 11054 6884 11056
rect 7376 11114 7436 11190
rect 7925 11248 9276 11250
rect 7925 11192 7930 11248
rect 7986 11192 9276 11248
rect 7925 11190 9276 11192
rect 9673 11250 9739 11253
rect 10726 11250 10732 11252
rect 9673 11248 10732 11250
rect 9673 11192 9678 11248
rect 9734 11192 10732 11248
rect 9673 11190 10732 11192
rect 7925 11187 7991 11190
rect 9673 11187 9739 11190
rect 10726 11188 10732 11190
rect 10796 11188 10802 11252
rect 10961 11248 11027 11253
rect 10961 11192 10966 11248
rect 11022 11192 11027 11248
rect 10961 11187 11027 11192
rect 11102 11250 11162 11462
rect 13261 11520 13971 11522
rect 13261 11464 13266 11520
rect 13322 11464 13910 11520
rect 13966 11464 13971 11520
rect 13261 11462 13971 11464
rect 13261 11459 13327 11462
rect 13905 11459 13971 11462
rect 14038 11460 14044 11524
rect 14108 11522 14114 11524
rect 14365 11522 14431 11525
rect 14825 11524 14891 11525
rect 14108 11520 14431 11522
rect 14108 11464 14370 11520
rect 14426 11464 14431 11520
rect 14108 11462 14431 11464
rect 14108 11460 14114 11462
rect 14365 11459 14431 11462
rect 14774 11460 14780 11524
rect 14844 11522 14891 11524
rect 14844 11520 14936 11522
rect 14886 11464 14936 11520
rect 14844 11462 14936 11464
rect 14844 11460 14891 11462
rect 14825 11459 14891 11460
rect 11946 11456 12262 11457
rect 11946 11392 11952 11456
rect 12016 11392 12032 11456
rect 12096 11392 12112 11456
rect 12176 11392 12192 11456
rect 12256 11392 12262 11456
rect 11946 11391 12262 11392
rect 16946 11456 17262 11457
rect 16946 11392 16952 11456
rect 17016 11392 17032 11456
rect 17096 11392 17112 11456
rect 17176 11392 17192 11456
rect 17256 11392 17262 11456
rect 16946 11391 17262 11392
rect 12433 11386 12499 11389
rect 13905 11386 13971 11389
rect 12433 11384 13971 11386
rect 12433 11328 12438 11384
rect 12494 11328 13910 11384
rect 13966 11328 13971 11384
rect 12433 11326 13971 11328
rect 12433 11323 12499 11326
rect 13905 11323 13971 11326
rect 14181 11386 14247 11389
rect 16246 11386 16252 11388
rect 14181 11384 16252 11386
rect 14181 11328 14186 11384
rect 14242 11328 16252 11384
rect 14181 11326 16252 11328
rect 14181 11323 14247 11326
rect 16246 11324 16252 11326
rect 16316 11324 16322 11388
rect 15837 11250 15903 11253
rect 11102 11248 15903 11250
rect 11102 11192 15842 11248
rect 15898 11192 15903 11248
rect 11102 11190 15903 11192
rect 16254 11250 16314 11324
rect 17769 11250 17835 11253
rect 16254 11248 17835 11250
rect 16254 11192 17774 11248
rect 17830 11192 17835 11248
rect 16254 11190 17835 11192
rect 15837 11187 15903 11190
rect 17769 11187 17835 11190
rect 17953 11250 18019 11253
rect 19200 11250 20000 11280
rect 17953 11248 20000 11250
rect 17953 11192 17958 11248
rect 18014 11192 20000 11248
rect 17953 11190 20000 11192
rect 17953 11187 18019 11190
rect 19200 11160 20000 11190
rect 12065 11114 12131 11117
rect 13813 11116 13879 11117
rect 13813 11114 13860 11116
rect 7376 11112 12131 11114
rect 7376 11056 12070 11112
rect 12126 11056 12131 11112
rect 7376 11054 12131 11056
rect 5073 11051 5139 11054
rect 12065 11051 12131 11054
rect 12436 11054 13692 11114
rect 13768 11112 13860 11114
rect 13768 11056 13818 11112
rect 13768 11054 13860 11056
rect 3182 10978 3188 10980
rect 3006 10918 3188 10978
rect 1117 10915 1183 10918
rect 3182 10916 3188 10918
rect 3252 10916 3258 10980
rect 3509 10978 3575 10981
rect 6177 10978 6243 10981
rect 6453 10978 6519 10981
rect 6913 10978 6979 10981
rect 3509 10976 5596 10978
rect 3509 10920 3514 10976
rect 3570 10920 5596 10976
rect 3509 10918 5596 10920
rect 3509 10915 3575 10918
rect 2606 10912 2922 10913
rect 2606 10848 2612 10912
rect 2676 10848 2692 10912
rect 2756 10848 2772 10912
rect 2836 10848 2852 10912
rect 2916 10848 2922 10912
rect 2606 10847 2922 10848
rect 3550 10780 3556 10844
rect 3620 10842 3626 10844
rect 4102 10842 4108 10844
rect 3620 10782 4108 10842
rect 3620 10780 3626 10782
rect 4102 10780 4108 10782
rect 4172 10780 4178 10844
rect 4286 10780 4292 10844
rect 4356 10842 4362 10844
rect 5390 10842 5396 10844
rect 4356 10782 5396 10842
rect 4356 10780 4362 10782
rect 5390 10780 5396 10782
rect 5460 10780 5466 10844
rect 5536 10842 5596 10918
rect 6177 10976 6519 10978
rect 6177 10920 6182 10976
rect 6238 10920 6458 10976
rect 6514 10920 6519 10976
rect 6177 10918 6519 10920
rect 6177 10915 6243 10918
rect 6453 10915 6519 10918
rect 6686 10976 6979 10978
rect 6686 10920 6918 10976
rect 6974 10920 6979 10976
rect 6686 10918 6979 10920
rect 6269 10842 6335 10845
rect 5536 10840 6335 10842
rect 5536 10784 6274 10840
rect 6330 10784 6335 10840
rect 5536 10782 6335 10784
rect 6269 10779 6335 10782
rect 2497 10706 2563 10709
rect 5441 10706 5507 10709
rect 6310 10706 6316 10708
rect 2497 10704 5507 10706
rect 2497 10648 2502 10704
rect 2558 10648 5446 10704
rect 5502 10648 5507 10704
rect 2497 10646 5507 10648
rect 2497 10643 2563 10646
rect 5441 10643 5507 10646
rect 5996 10646 6316 10706
rect 5996 10573 6056 10646
rect 6310 10644 6316 10646
rect 6380 10644 6386 10708
rect 6453 10706 6519 10709
rect 6686 10706 6746 10918
rect 6913 10915 6979 10918
rect 7281 10978 7347 10981
rect 7414 10978 7420 10980
rect 7281 10976 7420 10978
rect 7281 10920 7286 10976
rect 7342 10920 7420 10976
rect 7281 10918 7420 10920
rect 7281 10915 7347 10918
rect 7414 10916 7420 10918
rect 7484 10916 7490 10980
rect 9765 10978 9831 10981
rect 12436 10978 12496 11054
rect 9765 10976 12496 10978
rect 9765 10920 9770 10976
rect 9826 10920 12496 10976
rect 9765 10918 12496 10920
rect 13632 10978 13692 11054
rect 13813 11052 13860 11054
rect 13924 11052 13930 11116
rect 15878 11052 15884 11116
rect 15948 11114 15954 11116
rect 18137 11114 18203 11117
rect 15948 11112 18203 11114
rect 15948 11056 18142 11112
rect 18198 11056 18203 11112
rect 15948 11054 18203 11056
rect 15948 11052 15954 11054
rect 13813 11051 13879 11052
rect 18137 11051 18203 11054
rect 14590 10978 14596 10980
rect 13632 10918 14596 10978
rect 9765 10915 9831 10918
rect 14590 10916 14596 10918
rect 14660 10916 14666 10980
rect 15510 10916 15516 10980
rect 15580 10978 15586 10980
rect 17033 10978 17099 10981
rect 15580 10976 17099 10978
rect 15580 10920 17038 10976
rect 17094 10920 17099 10976
rect 15580 10918 17099 10920
rect 15580 10916 15586 10918
rect 17033 10915 17099 10918
rect 7606 10912 7922 10913
rect 7606 10848 7612 10912
rect 7676 10848 7692 10912
rect 7756 10848 7772 10912
rect 7836 10848 7852 10912
rect 7916 10848 7922 10912
rect 7606 10847 7922 10848
rect 12606 10912 12922 10913
rect 12606 10848 12612 10912
rect 12676 10848 12692 10912
rect 12756 10848 12772 10912
rect 12836 10848 12852 10912
rect 12916 10848 12922 10912
rect 12606 10847 12922 10848
rect 17606 10912 17922 10913
rect 17606 10848 17612 10912
rect 17676 10848 17692 10912
rect 17756 10848 17772 10912
rect 17836 10848 17852 10912
rect 17916 10848 17922 10912
rect 17606 10847 17922 10848
rect 6821 10842 6887 10845
rect 7414 10842 7420 10844
rect 6821 10840 7420 10842
rect 6821 10784 6826 10840
rect 6882 10784 7420 10840
rect 6821 10782 7420 10784
rect 6821 10779 6887 10782
rect 7414 10780 7420 10782
rect 7484 10780 7490 10844
rect 9949 10842 10015 10845
rect 8020 10840 10015 10842
rect 8020 10784 9954 10840
rect 10010 10784 10015 10840
rect 8020 10782 10015 10784
rect 7005 10706 7071 10709
rect 6453 10704 7071 10706
rect 6453 10648 6458 10704
rect 6514 10648 7010 10704
rect 7066 10648 7071 10704
rect 6453 10646 7071 10648
rect 6453 10643 6519 10646
rect 7005 10643 7071 10646
rect 7465 10706 7531 10709
rect 8020 10706 8080 10782
rect 9949 10779 10015 10782
rect 10726 10780 10732 10844
rect 10796 10842 10802 10844
rect 10961 10842 11027 10845
rect 10796 10840 11027 10842
rect 10796 10784 10966 10840
rect 11022 10784 11027 10840
rect 10796 10782 11027 10784
rect 10796 10780 10802 10782
rect 10961 10779 11027 10782
rect 11278 10780 11284 10844
rect 11348 10842 11354 10844
rect 12433 10842 12499 10845
rect 11348 10840 12499 10842
rect 11348 10784 12438 10840
rect 12494 10784 12499 10840
rect 11348 10782 12499 10784
rect 11348 10780 11354 10782
rect 12433 10779 12499 10782
rect 13261 10842 13327 10845
rect 14549 10842 14615 10845
rect 13261 10840 14615 10842
rect 13261 10784 13266 10840
rect 13322 10784 14554 10840
rect 14610 10784 14615 10840
rect 13261 10782 14615 10784
rect 13261 10779 13327 10782
rect 14549 10779 14615 10782
rect 14825 10842 14891 10845
rect 15285 10844 15351 10845
rect 15929 10844 15995 10845
rect 15285 10842 15332 10844
rect 14825 10840 15332 10842
rect 14825 10784 14830 10840
rect 14886 10784 15290 10840
rect 14825 10782 15332 10784
rect 14825 10779 14891 10782
rect 15285 10780 15332 10782
rect 15396 10780 15402 10844
rect 15878 10842 15884 10844
rect 15838 10782 15884 10842
rect 15948 10840 15995 10844
rect 15990 10784 15995 10840
rect 15878 10780 15884 10782
rect 15948 10780 15995 10784
rect 15285 10779 15351 10780
rect 15929 10779 15995 10780
rect 10961 10706 11027 10709
rect 11094 10706 11100 10708
rect 7465 10704 8080 10706
rect 7465 10648 7470 10704
rect 7526 10648 8080 10704
rect 7465 10646 8080 10648
rect 8158 10646 10840 10706
rect 7465 10643 7531 10646
rect 3049 10570 3115 10573
rect 3049 10568 4170 10570
rect 3049 10512 3054 10568
rect 3110 10512 4170 10568
rect 3049 10510 4170 10512
rect 3049 10507 3115 10510
rect 2773 10434 2839 10437
rect 3550 10434 3556 10436
rect 2773 10432 3556 10434
rect 2773 10376 2778 10432
rect 2834 10376 3556 10432
rect 2773 10374 3556 10376
rect 2773 10371 2839 10374
rect 3550 10372 3556 10374
rect 3620 10372 3626 10436
rect 3734 10372 3740 10436
rect 3804 10434 3810 10436
rect 3969 10434 4035 10437
rect 3804 10432 4035 10434
rect 3804 10376 3974 10432
rect 4030 10376 4035 10432
rect 3804 10374 4035 10376
rect 4110 10434 4170 10510
rect 5993 10568 6059 10573
rect 5993 10512 5998 10568
rect 6054 10512 6059 10568
rect 5993 10507 6059 10512
rect 6310 10508 6316 10572
rect 6380 10570 6386 10572
rect 6453 10570 6519 10573
rect 8158 10570 8218 10646
rect 6380 10568 6519 10570
rect 6380 10512 6458 10568
rect 6514 10512 6519 10568
rect 6380 10510 6519 10512
rect 6380 10508 6386 10510
rect 6453 10507 6519 10510
rect 6640 10510 8218 10570
rect 8569 10570 8635 10573
rect 9438 10570 9444 10572
rect 8569 10568 9444 10570
rect 8569 10512 8574 10568
rect 8630 10512 9444 10568
rect 8569 10510 9444 10512
rect 6640 10434 6700 10510
rect 8569 10507 8635 10510
rect 9438 10508 9444 10510
rect 9508 10508 9514 10572
rect 10780 10570 10840 10646
rect 10961 10704 11100 10706
rect 10961 10648 10966 10704
rect 11022 10648 11100 10704
rect 10961 10646 11100 10648
rect 10961 10643 11027 10646
rect 11094 10644 11100 10646
rect 11164 10644 11170 10708
rect 11513 10706 11579 10709
rect 17953 10706 18019 10709
rect 11513 10704 18019 10706
rect 11513 10648 11518 10704
rect 11574 10648 17958 10704
rect 18014 10648 18019 10704
rect 11513 10646 18019 10648
rect 11513 10643 11579 10646
rect 17953 10643 18019 10646
rect 11237 10570 11303 10573
rect 17493 10570 17559 10573
rect 10780 10568 11303 10570
rect 10780 10512 11242 10568
rect 11298 10512 11303 10568
rect 10780 10510 11303 10512
rect 11237 10507 11303 10510
rect 11424 10568 17559 10570
rect 11424 10512 17498 10568
rect 17554 10512 17559 10568
rect 11424 10510 17559 10512
rect 4110 10374 6700 10434
rect 7465 10434 7531 10437
rect 11424 10434 11484 10510
rect 17493 10507 17559 10510
rect 7465 10432 11484 10434
rect 7465 10376 7470 10432
rect 7526 10376 11484 10432
rect 7465 10374 11484 10376
rect 12709 10434 12775 10437
rect 15929 10434 15995 10437
rect 12709 10432 15995 10434
rect 12709 10376 12714 10432
rect 12770 10376 15934 10432
rect 15990 10376 15995 10432
rect 12709 10374 15995 10376
rect 3804 10372 3810 10374
rect 3969 10371 4035 10374
rect 7465 10371 7531 10374
rect 12709 10371 12775 10374
rect 15929 10371 15995 10374
rect 1946 10368 2262 10369
rect 1946 10304 1952 10368
rect 2016 10304 2032 10368
rect 2096 10304 2112 10368
rect 2176 10304 2192 10368
rect 2256 10304 2262 10368
rect 1946 10303 2262 10304
rect 6946 10368 7262 10369
rect 6946 10304 6952 10368
rect 7016 10304 7032 10368
rect 7096 10304 7112 10368
rect 7176 10304 7192 10368
rect 7256 10304 7262 10368
rect 6946 10303 7262 10304
rect 11946 10368 12262 10369
rect 11946 10304 11952 10368
rect 12016 10304 12032 10368
rect 12096 10304 12112 10368
rect 12176 10304 12192 10368
rect 12256 10304 12262 10368
rect 11946 10303 12262 10304
rect 16946 10368 17262 10369
rect 16946 10304 16952 10368
rect 17016 10304 17032 10368
rect 17096 10304 17112 10368
rect 17176 10304 17192 10368
rect 17256 10304 17262 10368
rect 16946 10303 17262 10304
rect 5758 10298 5764 10300
rect 3374 10238 5764 10298
rect 749 10162 815 10165
rect 3182 10162 3188 10164
rect 749 10160 3188 10162
rect 749 10104 754 10160
rect 810 10104 3188 10160
rect 749 10102 3188 10104
rect 749 10099 815 10102
rect 3182 10100 3188 10102
rect 3252 10100 3258 10164
rect 3374 10026 3434 10238
rect 5758 10236 5764 10238
rect 5828 10236 5834 10300
rect 7649 10298 7715 10301
rect 8201 10298 8267 10301
rect 9489 10300 9555 10301
rect 9438 10298 9444 10300
rect 7649 10296 8267 10298
rect 7649 10240 7654 10296
rect 7710 10240 8206 10296
rect 8262 10240 8267 10296
rect 7649 10238 8267 10240
rect 9398 10238 9444 10298
rect 9508 10296 9555 10300
rect 9550 10240 9555 10296
rect 7649 10235 7715 10238
rect 8201 10235 8267 10238
rect 9438 10236 9444 10238
rect 9508 10236 9555 10240
rect 9622 10236 9628 10300
rect 9692 10298 9698 10300
rect 10225 10298 10291 10301
rect 9692 10296 10291 10298
rect 9692 10240 10230 10296
rect 10286 10240 10291 10296
rect 9692 10238 10291 10240
rect 9692 10236 9698 10238
rect 9489 10235 9555 10236
rect 10225 10235 10291 10238
rect 10358 10236 10364 10300
rect 10428 10298 10434 10300
rect 11789 10298 11855 10301
rect 10428 10296 11855 10298
rect 10428 10240 11794 10296
rect 11850 10240 11855 10296
rect 10428 10238 11855 10240
rect 10428 10236 10434 10238
rect 11789 10235 11855 10238
rect 13486 10236 13492 10300
rect 13556 10298 13562 10300
rect 14457 10298 14523 10301
rect 13556 10296 14523 10298
rect 13556 10240 14462 10296
rect 14518 10240 14523 10296
rect 13556 10238 14523 10240
rect 13556 10236 13562 10238
rect 14457 10235 14523 10238
rect 15193 10298 15259 10301
rect 15837 10298 15903 10301
rect 15193 10296 15903 10298
rect 15193 10240 15198 10296
rect 15254 10240 15842 10296
rect 15898 10240 15903 10296
rect 15193 10238 15903 10240
rect 15193 10235 15259 10238
rect 15837 10235 15903 10238
rect 3509 10162 3575 10165
rect 3969 10162 4035 10165
rect 3509 10160 4035 10162
rect 3509 10104 3514 10160
rect 3570 10104 3974 10160
rect 4030 10104 4035 10160
rect 3509 10102 4035 10104
rect 3509 10099 3575 10102
rect 3969 10099 4035 10102
rect 4981 10162 5047 10165
rect 14181 10162 14247 10165
rect 4981 10160 14247 10162
rect 4981 10104 4986 10160
rect 5042 10104 14186 10160
rect 14242 10104 14247 10160
rect 4981 10102 14247 10104
rect 4981 10099 5047 10102
rect 14181 10099 14247 10102
rect 14549 10162 14615 10165
rect 15510 10162 15516 10164
rect 14549 10160 15516 10162
rect 14549 10104 14554 10160
rect 14610 10104 15516 10160
rect 14549 10102 15516 10104
rect 14549 10099 14615 10102
rect 15510 10100 15516 10102
rect 15580 10100 15586 10164
rect 16757 10162 16823 10165
rect 17769 10162 17835 10165
rect 16757 10160 17835 10162
rect 16757 10104 16762 10160
rect 16818 10104 17774 10160
rect 17830 10104 17835 10160
rect 16757 10102 17835 10104
rect 16757 10099 16823 10102
rect 17769 10099 17835 10102
rect 18137 10162 18203 10165
rect 19374 10162 19380 10164
rect 18137 10160 19380 10162
rect 18137 10104 18142 10160
rect 18198 10104 19380 10160
rect 18137 10102 19380 10104
rect 18137 10099 18203 10102
rect 19374 10100 19380 10102
rect 19444 10100 19450 10164
rect 2454 9966 3434 10026
rect 3601 10026 3667 10029
rect 4337 10028 4403 10029
rect 3601 10024 4216 10026
rect 3601 9968 3606 10024
rect 3662 9968 4216 10024
rect 3601 9966 4216 9968
rect 1025 9754 1091 9757
rect 1025 9752 1410 9754
rect 1025 9696 1030 9752
rect 1086 9696 1410 9752
rect 1025 9694 1410 9696
rect 1025 9691 1091 9694
rect 1350 9618 1410 9694
rect 2454 9621 2514 9966
rect 3601 9963 3667 9966
rect 2998 9828 3004 9892
rect 3068 9890 3074 9892
rect 3509 9890 3575 9893
rect 3068 9888 3575 9890
rect 3068 9832 3514 9888
rect 3570 9832 3575 9888
rect 3068 9830 3575 9832
rect 4156 9890 4216 9966
rect 4286 9964 4292 10028
rect 4356 10026 4403 10028
rect 4356 10024 4448 10026
rect 4398 9968 4448 10024
rect 4356 9966 4448 9968
rect 4356 9964 4403 9966
rect 5574 9964 5580 10028
rect 5644 10026 5650 10028
rect 6085 10026 6151 10029
rect 5644 10024 6151 10026
rect 5644 9968 6090 10024
rect 6146 9968 6151 10024
rect 5644 9966 6151 9968
rect 5644 9964 5650 9966
rect 4337 9963 4403 9964
rect 6085 9963 6151 9966
rect 6453 10026 6519 10029
rect 12249 10026 12315 10029
rect 17493 10026 17559 10029
rect 6453 10024 12315 10026
rect 6453 9968 6458 10024
rect 6514 9968 12254 10024
rect 12310 9968 12315 10024
rect 6453 9966 12315 9968
rect 6453 9963 6519 9966
rect 12249 9963 12315 9966
rect 12390 10024 17559 10026
rect 12390 9968 17498 10024
rect 17554 9968 17559 10024
rect 12390 9966 17559 9968
rect 8201 9890 8267 9893
rect 9489 9890 9555 9893
rect 4156 9830 7528 9890
rect 3068 9828 3074 9830
rect 3509 9827 3575 9830
rect 2606 9824 2922 9825
rect 2606 9760 2612 9824
rect 2676 9760 2692 9824
rect 2756 9760 2772 9824
rect 2836 9760 2852 9824
rect 2916 9760 2922 9824
rect 2606 9759 2922 9760
rect 3325 9754 3391 9757
rect 4337 9754 4403 9757
rect 3325 9752 4403 9754
rect 3325 9696 3330 9752
rect 3386 9696 4342 9752
rect 4398 9696 4403 9752
rect 3325 9694 4403 9696
rect 3325 9691 3391 9694
rect 4337 9691 4403 9694
rect 5257 9754 5323 9757
rect 5257 9752 6240 9754
rect 5257 9696 5262 9752
rect 5318 9696 6240 9752
rect 5257 9694 6240 9696
rect 5257 9691 5323 9694
rect 1350 9558 1778 9618
rect 1718 9484 1778 9558
rect 2405 9616 2514 9621
rect 2405 9560 2410 9616
rect 2466 9560 2514 9616
rect 2405 9558 2514 9560
rect 2865 9618 2931 9621
rect 3366 9618 3372 9620
rect 2865 9616 3372 9618
rect 2865 9560 2870 9616
rect 2926 9560 3372 9616
rect 2865 9558 3372 9560
rect 2405 9555 2471 9558
rect 2865 9555 2931 9558
rect 3366 9556 3372 9558
rect 3436 9556 3442 9620
rect 4797 9618 4863 9621
rect 5022 9618 5028 9620
rect 4797 9616 5028 9618
rect 4797 9560 4802 9616
rect 4858 9560 5028 9616
rect 4797 9558 5028 9560
rect 4797 9555 4863 9558
rect 5022 9556 5028 9558
rect 5092 9556 5098 9620
rect 6180 9618 6240 9694
rect 6310 9692 6316 9756
rect 6380 9754 6386 9756
rect 6453 9754 6519 9757
rect 6380 9752 6519 9754
rect 6380 9696 6458 9752
rect 6514 9696 6519 9752
rect 6380 9694 6519 9696
rect 6380 9692 6386 9694
rect 6453 9691 6519 9694
rect 6310 9618 6316 9620
rect 6180 9558 6316 9618
rect 6310 9556 6316 9558
rect 6380 9556 6386 9620
rect 7468 9618 7528 9830
rect 8201 9888 9555 9890
rect 8201 9832 8206 9888
rect 8262 9832 9494 9888
rect 9550 9832 9555 9888
rect 8201 9830 9555 9832
rect 8201 9827 8267 9830
rect 9489 9827 9555 9830
rect 11053 9890 11119 9893
rect 12390 9890 12450 9966
rect 17493 9963 17559 9966
rect 11053 9888 12450 9890
rect 11053 9832 11058 9888
rect 11114 9832 12450 9888
rect 11053 9830 12450 9832
rect 11053 9827 11119 9830
rect 13302 9828 13308 9892
rect 13372 9890 13378 9892
rect 13854 9890 13860 9892
rect 13372 9830 13860 9890
rect 13372 9828 13378 9830
rect 13854 9828 13860 9830
rect 13924 9828 13930 9892
rect 14181 9890 14247 9893
rect 15878 9890 15884 9892
rect 14181 9888 15884 9890
rect 14181 9832 14186 9888
rect 14242 9832 15884 9888
rect 14181 9830 15884 9832
rect 14181 9827 14247 9830
rect 15878 9828 15884 9830
rect 15948 9828 15954 9892
rect 16430 9828 16436 9892
rect 16500 9890 16506 9892
rect 17033 9890 17099 9893
rect 16500 9888 17099 9890
rect 16500 9832 17038 9888
rect 17094 9832 17099 9888
rect 16500 9830 17099 9832
rect 16500 9828 16506 9830
rect 17033 9827 17099 9830
rect 7606 9824 7922 9825
rect 7606 9760 7612 9824
rect 7676 9760 7692 9824
rect 7756 9760 7772 9824
rect 7836 9760 7852 9824
rect 7916 9760 7922 9824
rect 7606 9759 7922 9760
rect 12606 9824 12922 9825
rect 12606 9760 12612 9824
rect 12676 9760 12692 9824
rect 12756 9760 12772 9824
rect 12836 9760 12852 9824
rect 12916 9760 12922 9824
rect 12606 9759 12922 9760
rect 17606 9824 17922 9825
rect 17606 9760 17612 9824
rect 17676 9760 17692 9824
rect 17756 9760 17772 9824
rect 17836 9760 17852 9824
rect 17916 9760 17922 9824
rect 17606 9759 17922 9760
rect 9990 9754 9996 9756
rect 8020 9694 9996 9754
rect 8020 9618 8080 9694
rect 9990 9692 9996 9694
rect 10060 9692 10066 9756
rect 12157 9754 12223 9757
rect 12382 9754 12388 9756
rect 12157 9752 12388 9754
rect 12157 9696 12162 9752
rect 12218 9696 12388 9752
rect 12157 9694 12388 9696
rect 12157 9691 12223 9694
rect 12382 9692 12388 9694
rect 12452 9692 12458 9756
rect 13261 9754 13327 9757
rect 13486 9754 13492 9756
rect 13261 9752 13492 9754
rect 13261 9696 13266 9752
rect 13322 9696 13492 9752
rect 13261 9694 13492 9696
rect 13261 9691 13327 9694
rect 13486 9692 13492 9694
rect 13556 9692 13562 9756
rect 16062 9692 16068 9756
rect 16132 9754 16138 9756
rect 16481 9754 16547 9757
rect 16132 9752 16547 9754
rect 16132 9696 16486 9752
rect 16542 9696 16547 9752
rect 16132 9694 16547 9696
rect 16132 9692 16138 9694
rect 16481 9691 16547 9694
rect 18086 9692 18092 9756
rect 18156 9754 18162 9756
rect 18413 9754 18479 9757
rect 18156 9752 18479 9754
rect 18156 9696 18418 9752
rect 18474 9696 18479 9752
rect 18156 9694 18479 9696
rect 18156 9692 18162 9694
rect 18413 9691 18479 9694
rect 15101 9618 15167 9621
rect 7468 9558 8080 9618
rect 8204 9616 15167 9618
rect 8204 9560 15106 9616
rect 15162 9560 15167 9616
rect 8204 9558 15167 9560
rect 1710 9420 1716 9484
rect 1780 9482 1786 9484
rect 2037 9482 2103 9485
rect 1780 9480 2103 9482
rect 1780 9424 2042 9480
rect 2098 9424 2103 9480
rect 1780 9422 2103 9424
rect 1780 9420 1786 9422
rect 2037 9419 2103 9422
rect 2446 9420 2452 9484
rect 2516 9482 2522 9484
rect 2589 9482 2655 9485
rect 2516 9480 2655 9482
rect 2516 9424 2594 9480
rect 2650 9424 2655 9480
rect 2516 9422 2655 9424
rect 2516 9420 2522 9422
rect 2589 9419 2655 9422
rect 2957 9482 3023 9485
rect 3182 9482 3188 9484
rect 2957 9480 3188 9482
rect 2957 9424 2962 9480
rect 3018 9424 3188 9480
rect 2957 9422 3188 9424
rect 2957 9419 3023 9422
rect 3182 9420 3188 9422
rect 3252 9420 3258 9484
rect 3601 9482 3667 9485
rect 4889 9482 4955 9485
rect 3601 9480 4955 9482
rect 3601 9424 3606 9480
rect 3662 9424 4894 9480
rect 4950 9424 4955 9480
rect 3601 9422 4955 9424
rect 3601 9419 3667 9422
rect 4889 9419 4955 9422
rect 5165 9482 5231 9485
rect 5574 9482 5580 9484
rect 5165 9480 5580 9482
rect 5165 9424 5170 9480
rect 5226 9424 5580 9480
rect 5165 9422 5580 9424
rect 5165 9419 5231 9422
rect 5574 9420 5580 9422
rect 5644 9420 5650 9484
rect 5758 9420 5764 9484
rect 5828 9482 5834 9484
rect 8204 9482 8264 9558
rect 15101 9555 15167 9558
rect 16246 9556 16252 9620
rect 16316 9618 16322 9620
rect 16481 9618 16547 9621
rect 16798 9618 16804 9620
rect 16316 9616 16804 9618
rect 16316 9560 16486 9616
rect 16542 9560 16804 9616
rect 16316 9558 16804 9560
rect 16316 9556 16322 9558
rect 16481 9555 16547 9558
rect 16798 9556 16804 9558
rect 16868 9556 16874 9620
rect 9070 9482 9076 9484
rect 5828 9422 8264 9482
rect 8342 9422 9076 9482
rect 5828 9420 5834 9422
rect 3049 9346 3115 9349
rect 3182 9346 3188 9348
rect 3049 9344 3188 9346
rect 3049 9288 3054 9344
rect 3110 9288 3188 9344
rect 3049 9286 3188 9288
rect 3049 9283 3115 9286
rect 3182 9284 3188 9286
rect 3252 9284 3258 9348
rect 3325 9346 3391 9349
rect 3877 9346 3943 9349
rect 3325 9344 3943 9346
rect 3325 9288 3330 9344
rect 3386 9288 3882 9344
rect 3938 9288 3943 9344
rect 3325 9286 3943 9288
rect 3325 9283 3391 9286
rect 3877 9283 3943 9286
rect 4061 9346 4127 9349
rect 5022 9346 5028 9348
rect 4061 9344 5028 9346
rect 4061 9288 4066 9344
rect 4122 9288 5028 9344
rect 4061 9286 5028 9288
rect 4061 9283 4127 9286
rect 5022 9284 5028 9286
rect 5092 9284 5098 9348
rect 5206 9284 5212 9348
rect 5276 9346 5282 9348
rect 6361 9346 6427 9349
rect 5276 9344 6427 9346
rect 5276 9288 6366 9344
rect 6422 9288 6427 9344
rect 5276 9286 6427 9288
rect 5276 9284 5282 9286
rect 6361 9283 6427 9286
rect 7373 9346 7439 9349
rect 8342 9346 8402 9422
rect 9070 9420 9076 9422
rect 9140 9420 9146 9484
rect 9857 9482 9923 9485
rect 15561 9482 15627 9485
rect 16246 9482 16252 9484
rect 9857 9480 15627 9482
rect 9857 9424 9862 9480
rect 9918 9424 15566 9480
rect 15622 9424 15627 9480
rect 9857 9422 15627 9424
rect 9857 9419 9923 9422
rect 15561 9419 15627 9422
rect 15702 9422 16252 9482
rect 7373 9344 8402 9346
rect 7373 9288 7378 9344
rect 7434 9288 8402 9344
rect 7373 9286 8402 9288
rect 9029 9346 9095 9349
rect 14273 9348 14339 9349
rect 14457 9348 14523 9349
rect 14222 9346 14228 9348
rect 9029 9344 11852 9346
rect 9029 9288 9034 9344
rect 9090 9288 11852 9344
rect 9029 9286 11852 9288
rect 14182 9286 14228 9346
rect 14292 9344 14339 9348
rect 14334 9288 14339 9344
rect 7373 9283 7439 9286
rect 9029 9283 9095 9286
rect 1946 9280 2262 9281
rect 1946 9216 1952 9280
rect 2016 9216 2032 9280
rect 2096 9216 2112 9280
rect 2176 9216 2192 9280
rect 2256 9216 2262 9280
rect 1946 9215 2262 9216
rect 6946 9280 7262 9281
rect 6946 9216 6952 9280
rect 7016 9216 7032 9280
rect 7096 9216 7112 9280
rect 7176 9216 7192 9280
rect 7256 9216 7262 9280
rect 6946 9215 7262 9216
rect 4654 9210 4660 9212
rect 2730 9150 4660 9210
rect 749 9076 815 9077
rect 749 9074 796 9076
rect 704 9072 796 9074
rect 704 9016 754 9072
rect 704 9014 796 9016
rect 749 9012 796 9014
rect 860 9012 866 9076
rect 1577 9074 1643 9077
rect 2497 9074 2563 9077
rect 2730 9074 2790 9150
rect 4654 9148 4660 9150
rect 4724 9148 4730 9212
rect 5993 9210 6059 9213
rect 6310 9210 6316 9212
rect 5993 9208 6316 9210
rect 5993 9152 5998 9208
rect 6054 9152 6316 9208
rect 5993 9150 6316 9152
rect 5993 9147 6059 9150
rect 6310 9148 6316 9150
rect 6380 9148 6386 9212
rect 7373 9210 7439 9213
rect 8150 9210 8156 9212
rect 7373 9208 8156 9210
rect 7373 9152 7378 9208
rect 7434 9152 8156 9208
rect 7373 9150 8156 9152
rect 7373 9147 7439 9150
rect 8150 9148 8156 9150
rect 8220 9148 8226 9212
rect 10174 9148 10180 9212
rect 10244 9210 10250 9212
rect 10777 9210 10843 9213
rect 10244 9208 10843 9210
rect 10244 9152 10782 9208
rect 10838 9152 10843 9208
rect 10244 9150 10843 9152
rect 10244 9148 10250 9150
rect 10777 9147 10843 9150
rect 1577 9072 2790 9074
rect 1577 9016 1582 9072
rect 1638 9016 2502 9072
rect 2558 9016 2790 9072
rect 1577 9014 2790 9016
rect 2957 9074 3023 9077
rect 4102 9074 4108 9076
rect 2957 9072 4108 9074
rect 2957 9016 2962 9072
rect 3018 9016 4108 9072
rect 2957 9014 4108 9016
rect 749 9011 815 9012
rect 1577 9011 1643 9014
rect 2497 9011 2563 9014
rect 2957 9011 3023 9014
rect 4102 9012 4108 9014
rect 4172 9012 4178 9076
rect 8109 9074 8175 9077
rect 4524 9072 8175 9074
rect 4524 9016 8114 9072
rect 8170 9016 8175 9072
rect 4524 9014 8175 9016
rect 2129 8938 2195 8941
rect 4153 8938 4219 8941
rect 2129 8936 4219 8938
rect 2129 8880 2134 8936
rect 2190 8880 4158 8936
rect 4214 8880 4219 8936
rect 2129 8878 4219 8880
rect 2129 8875 2195 8878
rect 4153 8875 4219 8878
rect 0 8802 800 8832
rect 1945 8802 2011 8805
rect 0 8800 2011 8802
rect 0 8744 1950 8800
rect 2006 8744 2011 8800
rect 0 8742 2011 8744
rect 0 8712 800 8742
rect 1945 8739 2011 8742
rect 3417 8802 3483 8805
rect 3601 8802 3667 8805
rect 4524 8802 4584 9014
rect 8109 9011 8175 9014
rect 8886 9012 8892 9076
rect 8956 9074 8962 9076
rect 10501 9074 10567 9077
rect 8956 9072 10567 9074
rect 8956 9016 10506 9072
rect 10562 9016 10567 9072
rect 8956 9014 10567 9016
rect 8956 9012 8962 9014
rect 10501 9011 10567 9014
rect 10726 9012 10732 9076
rect 10796 9074 10802 9076
rect 10961 9074 11027 9077
rect 10796 9072 11027 9074
rect 10796 9016 10966 9072
rect 11022 9016 11027 9072
rect 10796 9014 11027 9016
rect 10796 9012 10802 9014
rect 10961 9011 11027 9014
rect 11278 9012 11284 9076
rect 11348 9074 11354 9076
rect 11605 9074 11671 9077
rect 11348 9072 11671 9074
rect 11348 9016 11610 9072
rect 11666 9016 11671 9072
rect 11348 9014 11671 9016
rect 11792 9074 11852 9286
rect 14222 9284 14228 9286
rect 14292 9284 14339 9288
rect 14406 9284 14412 9348
rect 14476 9346 14523 9348
rect 14476 9344 14568 9346
rect 14518 9288 14568 9344
rect 14476 9286 14568 9288
rect 14476 9284 14523 9286
rect 14273 9283 14339 9284
rect 14457 9283 14523 9284
rect 11946 9280 12262 9281
rect 11946 9216 11952 9280
rect 12016 9216 12032 9280
rect 12096 9216 12112 9280
rect 12176 9216 12192 9280
rect 12256 9216 12262 9280
rect 11946 9215 12262 9216
rect 15702 9210 15762 9422
rect 16246 9420 16252 9422
rect 16316 9482 16322 9484
rect 19149 9482 19215 9485
rect 16316 9480 19215 9482
rect 16316 9424 19154 9480
rect 19210 9424 19215 9480
rect 16316 9422 19215 9424
rect 16316 9420 16322 9422
rect 19149 9419 19215 9422
rect 16946 9280 17262 9281
rect 16946 9216 16952 9280
rect 17016 9216 17032 9280
rect 17096 9216 17112 9280
rect 17176 9216 17192 9280
rect 17256 9216 17262 9280
rect 16946 9215 17262 9216
rect 12390 9150 15762 9210
rect 12390 9074 12450 9150
rect 11792 9014 12450 9074
rect 12525 9074 12591 9077
rect 18137 9074 18203 9077
rect 12525 9072 18203 9074
rect 12525 9016 12530 9072
rect 12586 9016 18142 9072
rect 18198 9016 18203 9072
rect 12525 9014 18203 9016
rect 11348 9012 11354 9014
rect 11605 9011 11671 9014
rect 12525 9011 12591 9014
rect 18137 9011 18203 9014
rect 4654 8876 4660 8940
rect 4724 8938 4730 8940
rect 5349 8938 5415 8941
rect 4724 8936 5415 8938
rect 4724 8880 5354 8936
rect 5410 8880 5415 8936
rect 4724 8878 5415 8880
rect 4724 8876 4730 8878
rect 5349 8875 5415 8878
rect 6310 8876 6316 8940
rect 6380 8938 6386 8940
rect 7373 8938 7439 8941
rect 6380 8936 7439 8938
rect 6380 8880 7378 8936
rect 7434 8880 7439 8936
rect 6380 8878 7439 8880
rect 6380 8876 6386 8878
rect 7373 8875 7439 8878
rect 7649 8938 7715 8941
rect 9213 8938 9279 8941
rect 15653 8938 15719 8941
rect 18045 8938 18111 8941
rect 7649 8936 15719 8938
rect 7649 8880 7654 8936
rect 7710 8880 9218 8936
rect 9274 8880 15658 8936
rect 15714 8880 15719 8936
rect 7649 8878 15719 8880
rect 7649 8875 7715 8878
rect 9213 8875 9279 8878
rect 15653 8875 15719 8878
rect 15840 8936 18111 8938
rect 15840 8880 18050 8936
rect 18106 8880 18111 8936
rect 15840 8878 18111 8880
rect 3417 8800 3667 8802
rect 3417 8744 3422 8800
rect 3478 8744 3606 8800
rect 3662 8744 3667 8800
rect 3417 8742 3667 8744
rect 3417 8739 3483 8742
rect 3601 8739 3667 8742
rect 3880 8742 4584 8802
rect 5257 8802 5323 8805
rect 5257 8800 6608 8802
rect 5257 8744 5262 8800
rect 5318 8744 6608 8800
rect 5257 8742 6608 8744
rect 2606 8736 2922 8737
rect 2606 8672 2612 8736
rect 2676 8672 2692 8736
rect 2756 8672 2772 8736
rect 2836 8672 2852 8736
rect 2916 8672 2922 8736
rect 2606 8671 2922 8672
rect 1526 8604 1532 8668
rect 1596 8666 1602 8668
rect 2221 8666 2287 8669
rect 1596 8664 2287 8666
rect 1596 8608 2226 8664
rect 2282 8608 2287 8664
rect 1596 8606 2287 8608
rect 1596 8604 1602 8606
rect 2221 8603 2287 8606
rect 3880 8533 3940 8742
rect 5257 8739 5323 8742
rect 5390 8666 5396 8668
rect 4892 8606 5396 8666
rect 1342 8468 1348 8532
rect 1412 8530 1418 8532
rect 2589 8530 2655 8533
rect 1412 8528 2655 8530
rect 1412 8472 2594 8528
rect 2650 8472 2655 8528
rect 1412 8470 2655 8472
rect 1412 8468 1418 8470
rect 2589 8467 2655 8470
rect 2998 8468 3004 8532
rect 3068 8530 3074 8532
rect 3509 8530 3575 8533
rect 3068 8528 3575 8530
rect 3068 8472 3514 8528
rect 3570 8472 3575 8528
rect 3068 8470 3575 8472
rect 3068 8468 3074 8470
rect 3509 8467 3575 8470
rect 3877 8528 3943 8533
rect 3877 8472 3882 8528
rect 3938 8472 3943 8528
rect 3877 8467 3943 8472
rect 1301 8394 1367 8397
rect 3366 8394 3372 8396
rect 1301 8392 3372 8394
rect 1301 8336 1306 8392
rect 1362 8336 3372 8392
rect 1301 8334 3372 8336
rect 1301 8331 1367 8334
rect 3366 8332 3372 8334
rect 3436 8332 3442 8396
rect 3509 8394 3575 8397
rect 4892 8394 4952 8606
rect 5390 8604 5396 8606
rect 5460 8604 5466 8668
rect 6548 8666 6608 8742
rect 6678 8740 6684 8804
rect 6748 8802 6754 8804
rect 7373 8802 7439 8805
rect 6748 8800 7439 8802
rect 6748 8744 7378 8800
rect 7434 8744 7439 8800
rect 6748 8742 7439 8744
rect 6748 8740 6754 8742
rect 7373 8739 7439 8742
rect 8293 8802 8359 8805
rect 8886 8802 8892 8804
rect 8293 8800 8892 8802
rect 8293 8744 8298 8800
rect 8354 8744 8892 8800
rect 8293 8742 8892 8744
rect 8293 8739 8359 8742
rect 8886 8740 8892 8742
rect 8956 8740 8962 8804
rect 9765 8802 9831 8805
rect 12249 8802 12315 8805
rect 9765 8800 12315 8802
rect 9765 8744 9770 8800
rect 9826 8744 12254 8800
rect 12310 8744 12315 8800
rect 9765 8742 12315 8744
rect 9765 8739 9831 8742
rect 12249 8739 12315 8742
rect 14917 8802 14983 8805
rect 15840 8802 15900 8878
rect 18045 8875 18111 8878
rect 14917 8800 15900 8802
rect 14917 8744 14922 8800
rect 14978 8744 15900 8800
rect 14917 8742 15900 8744
rect 18413 8802 18479 8805
rect 19200 8802 20000 8832
rect 18413 8800 20000 8802
rect 18413 8744 18418 8800
rect 18474 8744 20000 8800
rect 18413 8742 20000 8744
rect 14917 8739 14983 8742
rect 18413 8739 18479 8742
rect 7606 8736 7922 8737
rect 7606 8672 7612 8736
rect 7676 8672 7692 8736
rect 7756 8672 7772 8736
rect 7836 8672 7852 8736
rect 7916 8672 7922 8736
rect 7606 8671 7922 8672
rect 12606 8736 12922 8737
rect 12606 8672 12612 8736
rect 12676 8672 12692 8736
rect 12756 8672 12772 8736
rect 12836 8672 12852 8736
rect 12916 8672 12922 8736
rect 12606 8671 12922 8672
rect 17606 8736 17922 8737
rect 17606 8672 17612 8736
rect 17676 8672 17692 8736
rect 17756 8672 17772 8736
rect 17836 8672 17852 8736
rect 17916 8672 17922 8736
rect 19200 8712 20000 8742
rect 17606 8671 17922 8672
rect 7005 8666 7071 8669
rect 6548 8664 7071 8666
rect 6548 8608 7010 8664
rect 7066 8608 7071 8664
rect 6548 8606 7071 8608
rect 7005 8603 7071 8606
rect 8385 8666 8451 8669
rect 10041 8666 10107 8669
rect 8385 8664 12450 8666
rect 8385 8608 8390 8664
rect 8446 8608 10046 8664
rect 10102 8608 12450 8664
rect 8385 8606 12450 8608
rect 8385 8603 8451 8606
rect 10041 8603 10107 8606
rect 5257 8530 5323 8533
rect 7281 8530 7347 8533
rect 9765 8530 9831 8533
rect 5257 8528 9831 8530
rect 5257 8472 5262 8528
rect 5318 8472 7286 8528
rect 7342 8472 9770 8528
rect 9826 8472 9831 8528
rect 5257 8470 9831 8472
rect 5257 8467 5323 8470
rect 7281 8467 7347 8470
rect 9765 8467 9831 8470
rect 9990 8468 9996 8532
rect 10060 8530 10066 8532
rect 10409 8530 10475 8533
rect 10060 8528 10475 8530
rect 10060 8472 10414 8528
rect 10470 8472 10475 8528
rect 10060 8470 10475 8472
rect 10060 8468 10066 8470
rect 10409 8467 10475 8470
rect 10777 8530 10843 8533
rect 11881 8530 11947 8533
rect 10777 8528 11947 8530
rect 10777 8472 10782 8528
rect 10838 8472 11886 8528
rect 11942 8472 11947 8528
rect 10777 8470 11947 8472
rect 12390 8530 12450 8606
rect 14549 8530 14615 8533
rect 18597 8530 18663 8533
rect 12390 8528 14615 8530
rect 12390 8472 14554 8528
rect 14610 8472 14615 8528
rect 12390 8470 14615 8472
rect 10777 8467 10843 8470
rect 11881 8467 11947 8470
rect 14549 8467 14615 8470
rect 16622 8528 18663 8530
rect 16622 8472 18602 8528
rect 18658 8472 18663 8528
rect 16622 8470 18663 8472
rect 3509 8392 4952 8394
rect 3509 8336 3514 8392
rect 3570 8336 4952 8392
rect 3509 8334 4952 8336
rect 5073 8394 5139 8397
rect 5390 8394 5396 8396
rect 5073 8392 5396 8394
rect 5073 8336 5078 8392
rect 5134 8336 5396 8392
rect 5073 8334 5396 8336
rect 3509 8331 3575 8334
rect 5073 8331 5139 8334
rect 5390 8332 5396 8334
rect 5460 8332 5466 8396
rect 5993 8394 6059 8397
rect 13302 8394 13308 8396
rect 5993 8392 13308 8394
rect 5993 8336 5998 8392
rect 6054 8336 13308 8392
rect 5993 8334 13308 8336
rect 5993 8331 6059 8334
rect 13302 8332 13308 8334
rect 13372 8394 13378 8396
rect 16622 8394 16682 8470
rect 18597 8467 18663 8470
rect 18873 8394 18939 8397
rect 13372 8334 16682 8394
rect 16760 8392 18939 8394
rect 16760 8336 18878 8392
rect 18934 8336 18939 8392
rect 16760 8334 18939 8336
rect 13372 8332 13378 8334
rect 4102 8196 4108 8260
rect 4172 8258 4178 8260
rect 4613 8258 4679 8261
rect 4172 8256 4679 8258
rect 4172 8200 4618 8256
rect 4674 8200 4679 8256
rect 4172 8198 4679 8200
rect 4172 8196 4178 8198
rect 4613 8195 4679 8198
rect 4889 8258 4955 8261
rect 6637 8260 6703 8261
rect 4889 8256 6562 8258
rect 4889 8200 4894 8256
rect 4950 8200 6562 8256
rect 4889 8198 6562 8200
rect 4889 8195 4955 8198
rect 1946 8192 2262 8193
rect 1946 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2262 8192
rect 1946 8127 2262 8128
rect 3049 8122 3115 8125
rect 3601 8122 3667 8125
rect 3049 8120 3667 8122
rect 3049 8064 3054 8120
rect 3110 8064 3606 8120
rect 3662 8064 3667 8120
rect 3049 8062 3667 8064
rect 3049 8059 3115 8062
rect 3601 8059 3667 8062
rect 3734 8060 3740 8124
rect 3804 8122 3810 8124
rect 3969 8122 4035 8125
rect 3804 8120 4035 8122
rect 3804 8064 3974 8120
rect 4030 8064 4035 8120
rect 3804 8062 4035 8064
rect 3804 8060 3810 8062
rect 3969 8059 4035 8062
rect 5257 8122 5323 8125
rect 5942 8122 5948 8124
rect 5257 8120 5948 8122
rect 5257 8064 5262 8120
rect 5318 8064 5948 8120
rect 5257 8062 5948 8064
rect 5257 8059 5323 8062
rect 5942 8060 5948 8062
rect 6012 8060 6018 8124
rect 6502 8122 6562 8198
rect 6637 8256 6684 8260
rect 6748 8258 6754 8260
rect 6637 8200 6642 8256
rect 6637 8196 6684 8200
rect 6748 8198 6794 8258
rect 6748 8196 6754 8198
rect 7414 8196 7420 8260
rect 7484 8258 7490 8260
rect 7557 8258 7623 8261
rect 7484 8256 7623 8258
rect 7484 8200 7562 8256
rect 7618 8200 7623 8256
rect 7484 8198 7623 8200
rect 7484 8196 7490 8198
rect 6637 8195 6703 8196
rect 7557 8195 7623 8198
rect 7925 8258 7991 8261
rect 8334 8258 8340 8260
rect 7925 8256 8340 8258
rect 7925 8200 7930 8256
rect 7986 8200 8340 8256
rect 7925 8198 8340 8200
rect 7925 8195 7991 8198
rect 8334 8196 8340 8198
rect 8404 8196 8410 8260
rect 9765 8258 9831 8261
rect 10726 8258 10732 8260
rect 9765 8256 10732 8258
rect 9765 8200 9770 8256
rect 9826 8200 10732 8256
rect 9765 8198 10732 8200
rect 9765 8195 9831 8198
rect 10726 8196 10732 8198
rect 10796 8196 10802 8260
rect 12985 8258 13051 8261
rect 13721 8258 13787 8261
rect 16760 8258 16820 8334
rect 18873 8331 18939 8334
rect 12985 8256 13787 8258
rect 12985 8200 12990 8256
rect 13046 8200 13726 8256
rect 13782 8200 13787 8256
rect 12985 8198 13787 8200
rect 12985 8195 13051 8198
rect 13721 8195 13787 8198
rect 13862 8198 16820 8258
rect 6946 8192 7262 8193
rect 6946 8128 6952 8192
rect 7016 8128 7032 8192
rect 7096 8128 7112 8192
rect 7176 8128 7192 8192
rect 7256 8128 7262 8192
rect 6946 8127 7262 8128
rect 11946 8192 12262 8193
rect 11946 8128 11952 8192
rect 12016 8128 12032 8192
rect 12096 8128 12112 8192
rect 12176 8128 12192 8192
rect 12256 8128 12262 8192
rect 11946 8127 12262 8128
rect 6729 8122 6795 8125
rect 6502 8120 6795 8122
rect 6502 8064 6734 8120
rect 6790 8064 6795 8120
rect 6502 8062 6795 8064
rect 6729 8059 6795 8062
rect 7557 8122 7623 8125
rect 9438 8122 9444 8124
rect 7557 8120 9444 8122
rect 7557 8064 7562 8120
rect 7618 8064 9444 8120
rect 7557 8062 9444 8064
rect 7557 8059 7623 8062
rect 9438 8060 9444 8062
rect 9508 8060 9514 8124
rect 9581 8122 9647 8125
rect 9949 8122 10015 8125
rect 9581 8120 10015 8122
rect 9581 8064 9586 8120
rect 9642 8064 9954 8120
rect 10010 8064 10015 8120
rect 9581 8062 10015 8064
rect 9581 8059 9647 8062
rect 9949 8059 10015 8062
rect 12617 8122 12683 8125
rect 13862 8122 13922 8198
rect 16946 8192 17262 8193
rect 16946 8128 16952 8192
rect 17016 8128 17032 8192
rect 17096 8128 17112 8192
rect 17176 8128 17192 8192
rect 17256 8128 17262 8192
rect 16946 8127 17262 8128
rect 12617 8120 13922 8122
rect 12617 8064 12622 8120
rect 12678 8064 13922 8120
rect 12617 8062 13922 8064
rect 12617 8059 12683 8062
rect 14590 8060 14596 8124
rect 14660 8122 14666 8124
rect 15101 8122 15167 8125
rect 14660 8120 15167 8122
rect 14660 8064 15106 8120
rect 15162 8064 15167 8120
rect 14660 8062 15167 8064
rect 14660 8060 14666 8062
rect 15101 8059 15167 8062
rect 3550 7924 3556 7988
rect 3620 7986 3626 7988
rect 7097 7986 7163 7989
rect 7741 7986 7807 7989
rect 8109 7988 8175 7989
rect 8109 7986 8156 7988
rect 3620 7926 5780 7986
rect 3620 7924 3626 7926
rect 3785 7850 3851 7853
rect 4654 7850 4660 7852
rect 3785 7848 4660 7850
rect 3785 7792 3790 7848
rect 3846 7792 4660 7848
rect 3785 7790 4660 7792
rect 3785 7787 3851 7790
rect 4654 7788 4660 7790
rect 4724 7788 4730 7852
rect 5720 7850 5780 7926
rect 7097 7984 7807 7986
rect 7097 7928 7102 7984
rect 7158 7928 7746 7984
rect 7802 7928 7807 7984
rect 7097 7926 7807 7928
rect 8064 7984 8156 7986
rect 8064 7928 8114 7984
rect 8064 7926 8156 7928
rect 7097 7923 7163 7926
rect 7741 7923 7807 7926
rect 8109 7924 8156 7926
rect 8220 7924 8226 7988
rect 8293 7986 8359 7989
rect 11329 7986 11395 7989
rect 13905 7986 13971 7989
rect 8293 7984 11395 7986
rect 8293 7928 8298 7984
rect 8354 7928 11334 7984
rect 11390 7928 11395 7984
rect 8293 7926 11395 7928
rect 8109 7923 8175 7924
rect 8293 7923 8359 7926
rect 11329 7923 11395 7926
rect 12252 7984 13971 7986
rect 12252 7928 13910 7984
rect 13966 7928 13971 7984
rect 12252 7926 13971 7928
rect 5720 7790 8080 7850
rect 5022 7652 5028 7716
rect 5092 7714 5098 7716
rect 7189 7714 7255 7717
rect 5092 7712 7255 7714
rect 5092 7656 7194 7712
rect 7250 7656 7255 7712
rect 5092 7654 7255 7656
rect 8020 7714 8080 7790
rect 8334 7788 8340 7852
rect 8404 7850 8410 7852
rect 12252 7850 12312 7926
rect 13905 7923 13971 7926
rect 15694 7924 15700 7988
rect 15764 7986 15770 7988
rect 16205 7986 16271 7989
rect 15764 7984 16271 7986
rect 15764 7928 16210 7984
rect 16266 7928 16271 7984
rect 15764 7926 16271 7928
rect 15764 7924 15770 7926
rect 16205 7923 16271 7926
rect 17033 7850 17099 7853
rect 17585 7850 17651 7853
rect 8404 7790 12312 7850
rect 12436 7848 17099 7850
rect 12436 7792 17038 7848
rect 17094 7792 17099 7848
rect 12436 7790 17099 7792
rect 8404 7788 8410 7790
rect 9489 7714 9555 7717
rect 8020 7712 9555 7714
rect 8020 7656 9494 7712
rect 9550 7656 9555 7712
rect 8020 7654 9555 7656
rect 5092 7652 5098 7654
rect 7189 7651 7255 7654
rect 9489 7651 9555 7654
rect 9673 7714 9739 7717
rect 11094 7714 11100 7716
rect 9673 7712 11100 7714
rect 9673 7656 9678 7712
rect 9734 7656 11100 7712
rect 9673 7654 11100 7656
rect 9673 7651 9739 7654
rect 11094 7652 11100 7654
rect 11164 7652 11170 7716
rect 11462 7652 11468 7716
rect 11532 7714 11538 7716
rect 11605 7714 11671 7717
rect 11532 7712 11671 7714
rect 11532 7656 11610 7712
rect 11666 7656 11671 7712
rect 11532 7654 11671 7656
rect 11532 7652 11538 7654
rect 11605 7651 11671 7654
rect 2606 7648 2922 7649
rect 2606 7584 2612 7648
rect 2676 7584 2692 7648
rect 2756 7584 2772 7648
rect 2836 7584 2852 7648
rect 2916 7584 2922 7648
rect 2606 7583 2922 7584
rect 7606 7648 7922 7649
rect 7606 7584 7612 7648
rect 7676 7584 7692 7648
rect 7756 7584 7772 7648
rect 7836 7584 7852 7648
rect 7916 7584 7922 7648
rect 7606 7583 7922 7584
rect 5942 7516 5948 7580
rect 6012 7578 6018 7580
rect 6453 7578 6519 7581
rect 12436 7578 12496 7790
rect 17033 7787 17099 7790
rect 17358 7848 17651 7850
rect 17358 7792 17590 7848
rect 17646 7792 17651 7848
rect 17358 7790 17651 7792
rect 14825 7714 14891 7717
rect 17358 7714 17418 7790
rect 17585 7787 17651 7790
rect 14825 7712 17418 7714
rect 14825 7656 14830 7712
rect 14886 7656 17418 7712
rect 14825 7654 17418 7656
rect 14825 7651 14891 7654
rect 12606 7648 12922 7649
rect 12606 7584 12612 7648
rect 12676 7584 12692 7648
rect 12756 7584 12772 7648
rect 12836 7584 12852 7648
rect 12916 7584 12922 7648
rect 12606 7583 12922 7584
rect 17606 7648 17922 7649
rect 17606 7584 17612 7648
rect 17676 7584 17692 7648
rect 17756 7584 17772 7648
rect 17836 7584 17852 7648
rect 17916 7584 17922 7648
rect 17606 7583 17922 7584
rect 6012 7576 6519 7578
rect 6012 7520 6458 7576
rect 6514 7520 6519 7576
rect 6012 7518 6519 7520
rect 6012 7516 6018 7518
rect 6453 7515 6519 7518
rect 8158 7518 12496 7578
rect 3969 7442 4035 7445
rect 5022 7442 5028 7444
rect 3969 7440 5028 7442
rect 3969 7384 3974 7440
rect 4030 7384 5028 7440
rect 3969 7382 5028 7384
rect 3969 7379 4035 7382
rect 5022 7380 5028 7382
rect 5092 7442 5098 7444
rect 8158 7442 8218 7518
rect 5092 7382 8218 7442
rect 5092 7380 5098 7382
rect 8334 7380 8340 7444
rect 8404 7442 8410 7444
rect 11973 7442 12039 7445
rect 8404 7440 12039 7442
rect 8404 7384 11978 7440
rect 12034 7384 12039 7440
rect 8404 7382 12039 7384
rect 8404 7380 8410 7382
rect 11973 7379 12039 7382
rect 841 7306 907 7309
rect 3550 7306 3556 7308
rect 841 7304 3556 7306
rect 841 7248 846 7304
rect 902 7248 3556 7304
rect 841 7246 3556 7248
rect 841 7243 907 7246
rect 3550 7244 3556 7246
rect 3620 7244 3626 7308
rect 4705 7306 4771 7309
rect 6126 7306 6132 7308
rect 4705 7304 6132 7306
rect 4705 7248 4710 7304
rect 4766 7248 6132 7304
rect 4705 7246 6132 7248
rect 4705 7243 4771 7246
rect 6126 7244 6132 7246
rect 6196 7306 6202 7308
rect 7557 7306 7623 7309
rect 6196 7304 7623 7306
rect 6196 7248 7562 7304
rect 7618 7248 7623 7304
rect 6196 7246 7623 7248
rect 6196 7244 6202 7246
rect 7557 7243 7623 7246
rect 10726 7244 10732 7308
rect 10796 7306 10802 7308
rect 17033 7306 17099 7309
rect 10796 7304 17099 7306
rect 10796 7248 17038 7304
rect 17094 7248 17099 7304
rect 10796 7246 17099 7248
rect 10796 7244 10802 7246
rect 17033 7243 17099 7246
rect 1761 7172 1827 7173
rect 1710 7170 1716 7172
rect 1670 7110 1716 7170
rect 1780 7168 1827 7172
rect 1822 7112 1827 7168
rect 1710 7108 1716 7110
rect 1780 7108 1827 7112
rect 1761 7107 1827 7108
rect 8293 7170 8359 7173
rect 9305 7170 9371 7173
rect 8293 7168 9371 7170
rect 8293 7112 8298 7168
rect 8354 7112 9310 7168
rect 9366 7112 9371 7168
rect 8293 7110 9371 7112
rect 8293 7107 8359 7110
rect 9305 7107 9371 7110
rect 10358 7108 10364 7172
rect 10428 7170 10434 7172
rect 11605 7170 11671 7173
rect 10428 7168 11671 7170
rect 10428 7112 11610 7168
rect 11666 7112 11671 7168
rect 10428 7110 11671 7112
rect 10428 7108 10434 7110
rect 11605 7107 11671 7110
rect 12382 7108 12388 7172
rect 12452 7170 12458 7172
rect 13445 7170 13511 7173
rect 12452 7168 13511 7170
rect 12452 7112 13450 7168
rect 13506 7112 13511 7168
rect 12452 7110 13511 7112
rect 12452 7108 12458 7110
rect 13445 7107 13511 7110
rect 14365 7170 14431 7173
rect 14733 7170 14799 7173
rect 14365 7168 14799 7170
rect 14365 7112 14370 7168
rect 14426 7112 14738 7168
rect 14794 7112 14799 7168
rect 14365 7110 14799 7112
rect 14365 7107 14431 7110
rect 14733 7107 14799 7110
rect 1946 7104 2262 7105
rect 1946 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2262 7104
rect 1946 7039 2262 7040
rect 6946 7104 7262 7105
rect 6946 7040 6952 7104
rect 7016 7040 7032 7104
rect 7096 7040 7112 7104
rect 7176 7040 7192 7104
rect 7256 7040 7262 7104
rect 6946 7039 7262 7040
rect 11946 7104 12262 7105
rect 11946 7040 11952 7104
rect 12016 7040 12032 7104
rect 12096 7040 12112 7104
rect 12176 7040 12192 7104
rect 12256 7040 12262 7104
rect 11946 7039 12262 7040
rect 16946 7104 17262 7105
rect 16946 7040 16952 7104
rect 17016 7040 17032 7104
rect 17096 7040 17112 7104
rect 17176 7040 17192 7104
rect 17256 7040 17262 7104
rect 16946 7039 17262 7040
rect 3877 7036 3943 7037
rect 3877 7032 3924 7036
rect 3988 7034 3994 7036
rect 3877 6976 3882 7032
rect 3877 6972 3924 6976
rect 3988 6974 4034 7034
rect 3988 6972 3994 6974
rect 9438 6972 9444 7036
rect 9508 7034 9514 7036
rect 10777 7034 10843 7037
rect 11053 7036 11119 7037
rect 11053 7034 11100 7036
rect 9508 7032 10843 7034
rect 9508 6976 10782 7032
rect 10838 6976 10843 7032
rect 9508 6974 10843 6976
rect 11008 7032 11100 7034
rect 11008 6976 11058 7032
rect 11008 6974 11100 6976
rect 9508 6972 9514 6974
rect 3877 6971 3943 6972
rect 10777 6971 10843 6974
rect 11053 6972 11100 6974
rect 11164 6972 11170 7036
rect 15377 7034 15443 7037
rect 12436 7032 15443 7034
rect 12436 6976 15382 7032
rect 15438 6976 15443 7032
rect 12436 6974 15443 6976
rect 11053 6971 11119 6972
rect 381 6898 447 6901
rect 381 6896 3066 6898
rect 381 6840 386 6896
rect 442 6840 3066 6896
rect 381 6838 3066 6840
rect 381 6835 447 6838
rect 2221 6762 2287 6765
rect 2405 6762 2471 6765
rect 2221 6760 2471 6762
rect 2221 6704 2226 6760
rect 2282 6704 2410 6760
rect 2466 6704 2471 6760
rect 2221 6702 2471 6704
rect 2221 6699 2287 6702
rect 2405 6699 2471 6702
rect 3006 6626 3066 6838
rect 3366 6836 3372 6900
rect 3436 6898 3442 6900
rect 4061 6898 4127 6901
rect 3436 6896 4127 6898
rect 3436 6840 4066 6896
rect 4122 6840 4127 6896
rect 3436 6838 4127 6840
rect 3436 6836 3442 6838
rect 4061 6835 4127 6838
rect 5717 6898 5783 6901
rect 12436 6898 12496 6974
rect 15377 6971 15443 6974
rect 5717 6896 12496 6898
rect 5717 6840 5722 6896
rect 5778 6840 12496 6896
rect 5717 6838 12496 6840
rect 12617 6898 12683 6901
rect 13118 6898 13124 6900
rect 12617 6896 13124 6898
rect 12617 6840 12622 6896
rect 12678 6840 13124 6896
rect 12617 6838 13124 6840
rect 5717 6835 5783 6838
rect 12617 6835 12683 6838
rect 13118 6836 13124 6838
rect 13188 6836 13194 6900
rect 17493 6898 17559 6901
rect 14966 6896 17559 6898
rect 14966 6840 17498 6896
rect 17554 6840 17559 6896
rect 14966 6838 17559 6840
rect 6085 6762 6151 6765
rect 6269 6762 6335 6765
rect 6085 6760 6335 6762
rect 6085 6704 6090 6760
rect 6146 6704 6274 6760
rect 6330 6704 6335 6760
rect 6085 6702 6335 6704
rect 6085 6699 6151 6702
rect 6269 6699 6335 6702
rect 6494 6700 6500 6764
rect 6564 6762 6570 6764
rect 6637 6762 6703 6765
rect 6564 6760 6703 6762
rect 6564 6704 6642 6760
rect 6698 6704 6703 6760
rect 6564 6702 6703 6704
rect 6564 6700 6570 6702
rect 6637 6699 6703 6702
rect 7557 6762 7623 6765
rect 9029 6762 9095 6765
rect 7557 6760 9095 6762
rect 7557 6704 7562 6760
rect 7618 6704 9034 6760
rect 9090 6704 9095 6760
rect 7557 6702 9095 6704
rect 7557 6699 7623 6702
rect 9029 6699 9095 6702
rect 9581 6762 9647 6765
rect 14966 6762 15026 6838
rect 17493 6835 17559 6838
rect 9581 6760 15026 6762
rect 9581 6704 9586 6760
rect 9642 6704 15026 6760
rect 9581 6702 15026 6704
rect 15377 6762 15443 6765
rect 15694 6762 15700 6764
rect 15377 6760 15700 6762
rect 15377 6704 15382 6760
rect 15438 6704 15700 6760
rect 15377 6702 15700 6704
rect 9581 6699 9647 6702
rect 15377 6699 15443 6702
rect 15694 6700 15700 6702
rect 15764 6700 15770 6764
rect 4429 6626 4495 6629
rect 3006 6624 4495 6626
rect 3006 6568 4434 6624
rect 4490 6568 4495 6624
rect 3006 6566 4495 6568
rect 4429 6563 4495 6566
rect 4889 6626 4955 6629
rect 7373 6626 7439 6629
rect 4889 6624 7439 6626
rect 4889 6568 4894 6624
rect 4950 6568 7378 6624
rect 7434 6568 7439 6624
rect 4889 6566 7439 6568
rect 4889 6563 4955 6566
rect 7373 6563 7439 6566
rect 8937 6626 9003 6629
rect 9857 6626 9923 6629
rect 8937 6624 9923 6626
rect 8937 6568 8942 6624
rect 8998 6568 9862 6624
rect 9918 6568 9923 6624
rect 8937 6566 9923 6568
rect 8937 6563 9003 6566
rect 9857 6563 9923 6566
rect 13629 6626 13695 6629
rect 16205 6626 16271 6629
rect 13629 6624 16271 6626
rect 13629 6568 13634 6624
rect 13690 6568 16210 6624
rect 16266 6568 16271 6624
rect 13629 6566 16271 6568
rect 13629 6563 13695 6566
rect 16205 6563 16271 6566
rect 2606 6560 2922 6561
rect 2606 6496 2612 6560
rect 2676 6496 2692 6560
rect 2756 6496 2772 6560
rect 2836 6496 2852 6560
rect 2916 6496 2922 6560
rect 2606 6495 2922 6496
rect 7606 6560 7922 6561
rect 7606 6496 7612 6560
rect 7676 6496 7692 6560
rect 7756 6496 7772 6560
rect 7836 6496 7852 6560
rect 7916 6496 7922 6560
rect 7606 6495 7922 6496
rect 12606 6560 12922 6561
rect 12606 6496 12612 6560
rect 12676 6496 12692 6560
rect 12756 6496 12772 6560
rect 12836 6496 12852 6560
rect 12916 6496 12922 6560
rect 12606 6495 12922 6496
rect 17606 6560 17922 6561
rect 17606 6496 17612 6560
rect 17676 6496 17692 6560
rect 17756 6496 17772 6560
rect 17836 6496 17852 6560
rect 17916 6496 17922 6560
rect 17606 6495 17922 6496
rect 1526 6428 1532 6492
rect 1596 6490 1602 6492
rect 3325 6490 3391 6493
rect 7281 6490 7347 6493
rect 9581 6490 9647 6493
rect 1596 6430 1778 6490
rect 1596 6428 1602 6430
rect 0 6354 800 6384
rect 1485 6354 1551 6357
rect 0 6352 1551 6354
rect 0 6296 1490 6352
rect 1546 6296 1551 6352
rect 0 6294 1551 6296
rect 1718 6354 1778 6430
rect 3325 6488 7347 6490
rect 3325 6432 3330 6488
rect 3386 6432 7286 6488
rect 7342 6432 7347 6488
rect 3325 6430 7347 6432
rect 3325 6427 3391 6430
rect 7281 6427 7347 6430
rect 8020 6488 9647 6490
rect 8020 6432 9586 6488
rect 9642 6432 9647 6488
rect 8020 6430 9647 6432
rect 4153 6354 4219 6357
rect 8020 6354 8080 6430
rect 9581 6427 9647 6430
rect 9949 6490 10015 6493
rect 10174 6490 10180 6492
rect 9949 6488 10180 6490
rect 9949 6432 9954 6488
rect 10010 6432 10180 6488
rect 9949 6430 10180 6432
rect 9949 6427 10015 6430
rect 10174 6428 10180 6430
rect 10244 6428 10250 6492
rect 13670 6428 13676 6492
rect 13740 6490 13746 6492
rect 15694 6490 15700 6492
rect 13740 6430 15700 6490
rect 13740 6428 13746 6430
rect 15694 6428 15700 6430
rect 15764 6490 15770 6492
rect 16205 6490 16271 6493
rect 15764 6488 16271 6490
rect 15764 6432 16210 6488
rect 16266 6432 16271 6488
rect 15764 6430 16271 6432
rect 15764 6428 15770 6430
rect 16205 6427 16271 6430
rect 1718 6294 3572 6354
rect 0 6264 800 6294
rect 1485 6291 1551 6294
rect 3512 6221 3572 6294
rect 4153 6352 8080 6354
rect 4153 6296 4158 6352
rect 4214 6296 8080 6352
rect 4153 6294 8080 6296
rect 4153 6291 4219 6294
rect 8150 6292 8156 6356
rect 8220 6354 8226 6356
rect 9673 6354 9739 6357
rect 8220 6352 9739 6354
rect 8220 6296 9678 6352
rect 9734 6296 9739 6352
rect 8220 6294 9739 6296
rect 8220 6292 8226 6294
rect 9673 6291 9739 6294
rect 10358 6292 10364 6356
rect 10428 6354 10434 6356
rect 16021 6354 16087 6357
rect 10428 6352 16087 6354
rect 10428 6296 16026 6352
rect 16082 6296 16087 6352
rect 10428 6294 16087 6296
rect 10428 6292 10434 6294
rect 16021 6291 16087 6294
rect 18413 6354 18479 6357
rect 19200 6354 20000 6384
rect 18413 6352 20000 6354
rect 18413 6296 18418 6352
rect 18474 6296 20000 6352
rect 18413 6294 20000 6296
rect 18413 6291 18479 6294
rect 19200 6264 20000 6294
rect 2221 6218 2287 6221
rect 2221 6216 2790 6218
rect 2221 6160 2226 6216
rect 2282 6160 2790 6216
rect 2221 6158 2790 6160
rect 2221 6155 2287 6158
rect 2730 6082 2790 6158
rect 3509 6216 3575 6221
rect 3509 6160 3514 6216
rect 3570 6160 3575 6216
rect 3509 6155 3575 6160
rect 3969 6218 4035 6221
rect 4286 6218 4292 6220
rect 3969 6216 4292 6218
rect 3969 6160 3974 6216
rect 4030 6160 4292 6216
rect 3969 6158 4292 6160
rect 3969 6155 4035 6158
rect 4286 6156 4292 6158
rect 4356 6156 4362 6220
rect 4654 6156 4660 6220
rect 4724 6218 4730 6220
rect 4889 6218 4955 6221
rect 4724 6216 4955 6218
rect 4724 6160 4894 6216
rect 4950 6160 4955 6216
rect 4724 6158 4955 6160
rect 4724 6156 4730 6158
rect 4889 6155 4955 6158
rect 6269 6218 6335 6221
rect 6494 6218 6500 6220
rect 6269 6216 6500 6218
rect 6269 6160 6274 6216
rect 6330 6160 6500 6216
rect 6269 6158 6500 6160
rect 6269 6155 6335 6158
rect 6494 6156 6500 6158
rect 6564 6156 6570 6220
rect 6637 6218 6703 6221
rect 16757 6218 16823 6221
rect 6637 6216 16823 6218
rect 6637 6160 6642 6216
rect 6698 6160 16762 6216
rect 16818 6160 16823 6216
rect 6637 6158 16823 6160
rect 6637 6155 6703 6158
rect 16757 6155 16823 6158
rect 8017 6082 8083 6085
rect 11462 6082 11468 6084
rect 2730 6022 6792 6082
rect 1946 6016 2262 6017
rect 1946 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2262 6016
rect 1946 5951 2262 5952
rect 4061 5948 4127 5949
rect 4061 5946 4108 5948
rect 4016 5944 4108 5946
rect 4016 5888 4066 5944
rect 4016 5886 4108 5888
rect 4061 5884 4108 5886
rect 4172 5884 4178 5948
rect 5809 5946 5875 5949
rect 5942 5946 5948 5948
rect 5809 5944 5948 5946
rect 5809 5888 5814 5944
rect 5870 5888 5948 5944
rect 5809 5886 5948 5888
rect 4061 5883 4127 5884
rect 5809 5883 5875 5886
rect 5942 5884 5948 5886
rect 6012 5884 6018 5948
rect 3877 5810 3943 5813
rect 4838 5810 4844 5812
rect 3877 5808 4844 5810
rect 3877 5752 3882 5808
rect 3938 5752 4844 5808
rect 3877 5750 4844 5752
rect 3877 5747 3943 5750
rect 4838 5748 4844 5750
rect 4908 5748 4914 5812
rect 5758 5748 5764 5812
rect 5828 5810 5834 5812
rect 6453 5810 6519 5813
rect 5828 5808 6519 5810
rect 5828 5752 6458 5808
rect 6514 5752 6519 5808
rect 5828 5750 6519 5752
rect 6732 5810 6792 6022
rect 8017 6080 11468 6082
rect 8017 6024 8022 6080
rect 8078 6024 11468 6080
rect 8017 6022 11468 6024
rect 8017 6019 8083 6022
rect 11462 6020 11468 6022
rect 11532 6020 11538 6084
rect 12709 6082 12775 6085
rect 16481 6082 16547 6085
rect 12709 6080 16547 6082
rect 12709 6024 12714 6080
rect 12770 6024 16486 6080
rect 16542 6024 16547 6080
rect 12709 6022 16547 6024
rect 12709 6019 12775 6022
rect 16481 6019 16547 6022
rect 6946 6016 7262 6017
rect 6946 5952 6952 6016
rect 7016 5952 7032 6016
rect 7096 5952 7112 6016
rect 7176 5952 7192 6016
rect 7256 5952 7262 6016
rect 6946 5951 7262 5952
rect 11946 6016 12262 6017
rect 11946 5952 11952 6016
rect 12016 5952 12032 6016
rect 12096 5952 12112 6016
rect 12176 5952 12192 6016
rect 12256 5952 12262 6016
rect 11946 5951 12262 5952
rect 16946 6016 17262 6017
rect 16946 5952 16952 6016
rect 17016 5952 17032 6016
rect 17096 5952 17112 6016
rect 17176 5952 17192 6016
rect 17256 5952 17262 6016
rect 16946 5951 17262 5952
rect 7649 5946 7715 5949
rect 8150 5946 8156 5948
rect 7649 5944 8156 5946
rect 7649 5888 7654 5944
rect 7710 5888 8156 5944
rect 7649 5886 8156 5888
rect 7649 5883 7715 5886
rect 8150 5884 8156 5886
rect 8220 5884 8226 5948
rect 8937 5946 9003 5949
rect 9806 5946 9812 5948
rect 8937 5944 9812 5946
rect 8937 5888 8942 5944
rect 8998 5888 9812 5944
rect 8937 5886 9812 5888
rect 8937 5883 9003 5886
rect 9806 5884 9812 5886
rect 9876 5884 9882 5948
rect 12433 5946 12499 5949
rect 16573 5946 16639 5949
rect 12433 5944 16639 5946
rect 12433 5888 12438 5944
rect 12494 5888 16578 5944
rect 16634 5888 16639 5944
rect 12433 5886 16639 5888
rect 12433 5883 12499 5886
rect 16573 5883 16639 5886
rect 7005 5810 7071 5813
rect 9489 5810 9555 5813
rect 6732 5808 9555 5810
rect 6732 5752 7010 5808
rect 7066 5752 9494 5808
rect 9550 5752 9555 5808
rect 6732 5750 9555 5752
rect 5828 5748 5834 5750
rect 6453 5747 6519 5750
rect 7005 5747 7071 5750
rect 9489 5747 9555 5750
rect 10726 5748 10732 5812
rect 10796 5810 10802 5812
rect 18086 5810 18092 5812
rect 10796 5750 18092 5810
rect 10796 5748 10802 5750
rect 18086 5748 18092 5750
rect 18156 5748 18162 5812
rect 790 5612 796 5676
rect 860 5674 866 5676
rect 7097 5674 7163 5677
rect 14181 5674 14247 5677
rect 18270 5674 18276 5676
rect 860 5614 6930 5674
rect 860 5612 866 5614
rect 3509 5538 3575 5541
rect 6729 5538 6795 5541
rect 3509 5536 6795 5538
rect 3509 5480 3514 5536
rect 3570 5480 6734 5536
rect 6790 5480 6795 5536
rect 3509 5478 6795 5480
rect 6870 5538 6930 5614
rect 7097 5672 14247 5674
rect 7097 5616 7102 5672
rect 7158 5616 14186 5672
rect 14242 5616 14247 5672
rect 7097 5614 14247 5616
rect 7097 5611 7163 5614
rect 14181 5611 14247 5614
rect 16576 5614 18276 5674
rect 7281 5538 7347 5541
rect 6870 5536 7347 5538
rect 6870 5480 7286 5536
rect 7342 5480 7347 5536
rect 6870 5478 7347 5480
rect 3509 5475 3575 5478
rect 6729 5475 6795 5478
rect 7281 5475 7347 5478
rect 9121 5538 9187 5541
rect 9990 5538 9996 5540
rect 9121 5536 9996 5538
rect 9121 5480 9126 5536
rect 9182 5480 9996 5536
rect 9121 5478 9996 5480
rect 9121 5475 9187 5478
rect 9990 5476 9996 5478
rect 10060 5476 10066 5540
rect 10869 5536 10935 5541
rect 10869 5480 10874 5536
rect 10930 5480 10935 5536
rect 10869 5475 10935 5480
rect 11278 5476 11284 5540
rect 11348 5538 11354 5540
rect 11789 5538 11855 5541
rect 11348 5536 11855 5538
rect 11348 5480 11794 5536
rect 11850 5480 11855 5536
rect 11348 5478 11855 5480
rect 11348 5476 11354 5478
rect 11789 5475 11855 5478
rect 15929 5538 15995 5541
rect 16576 5538 16636 5614
rect 18270 5612 18276 5614
rect 18340 5612 18346 5676
rect 15929 5536 16636 5538
rect 15929 5480 15934 5536
rect 15990 5480 16636 5536
rect 15929 5478 16636 5480
rect 18321 5538 18387 5541
rect 18454 5538 18460 5540
rect 18321 5536 18460 5538
rect 18321 5480 18326 5536
rect 18382 5480 18460 5536
rect 18321 5478 18460 5480
rect 15929 5475 15995 5478
rect 18321 5475 18387 5478
rect 18454 5476 18460 5478
rect 18524 5476 18530 5540
rect 2606 5472 2922 5473
rect 2606 5408 2612 5472
rect 2676 5408 2692 5472
rect 2756 5408 2772 5472
rect 2836 5408 2852 5472
rect 2916 5408 2922 5472
rect 2606 5407 2922 5408
rect 7606 5472 7922 5473
rect 7606 5408 7612 5472
rect 7676 5408 7692 5472
rect 7756 5408 7772 5472
rect 7836 5408 7852 5472
rect 7916 5408 7922 5472
rect 7606 5407 7922 5408
rect 3969 5402 4035 5405
rect 7465 5402 7531 5405
rect 3969 5400 7531 5402
rect 3969 5344 3974 5400
rect 4030 5344 7470 5400
rect 7526 5344 7531 5400
rect 3969 5342 7531 5344
rect 3969 5339 4035 5342
rect 7465 5339 7531 5342
rect 8385 5402 8451 5405
rect 10872 5402 10932 5475
rect 12606 5472 12922 5473
rect 12606 5408 12612 5472
rect 12676 5408 12692 5472
rect 12756 5408 12772 5472
rect 12836 5408 12852 5472
rect 12916 5408 12922 5472
rect 12606 5407 12922 5408
rect 17606 5472 17922 5473
rect 17606 5408 17612 5472
rect 17676 5408 17692 5472
rect 17756 5408 17772 5472
rect 17836 5408 17852 5472
rect 17916 5408 17922 5472
rect 17606 5407 17922 5408
rect 11278 5402 11284 5404
rect 8385 5400 11284 5402
rect 8385 5344 8390 5400
rect 8446 5344 11284 5400
rect 8385 5342 11284 5344
rect 8385 5339 8451 5342
rect 11278 5340 11284 5342
rect 11348 5340 11354 5404
rect 12249 5402 12315 5405
rect 12382 5402 12388 5404
rect 12249 5400 12388 5402
rect 12249 5344 12254 5400
rect 12310 5344 12388 5400
rect 12249 5342 12388 5344
rect 12249 5339 12315 5342
rect 12382 5340 12388 5342
rect 12452 5340 12458 5404
rect 3049 5268 3115 5269
rect 2998 5266 3004 5268
rect 2958 5206 3004 5266
rect 3068 5264 3115 5268
rect 3110 5208 3115 5264
rect 2998 5204 3004 5206
rect 3068 5204 3115 5208
rect 5574 5204 5580 5268
rect 5644 5266 5650 5268
rect 5717 5266 5783 5269
rect 5644 5264 5783 5266
rect 5644 5208 5722 5264
rect 5778 5208 5783 5264
rect 5644 5206 5783 5208
rect 5644 5204 5650 5206
rect 3049 5203 3115 5204
rect 5717 5203 5783 5206
rect 6678 5204 6684 5268
rect 6748 5266 6754 5268
rect 8845 5266 8911 5269
rect 6748 5264 8911 5266
rect 6748 5208 8850 5264
rect 8906 5208 8911 5264
rect 6748 5206 8911 5208
rect 6748 5204 6754 5206
rect 8845 5203 8911 5206
rect 9070 5204 9076 5268
rect 9140 5266 9146 5268
rect 11513 5266 11579 5269
rect 13302 5266 13308 5268
rect 9140 5206 11070 5266
rect 9140 5204 9146 5206
rect 974 5068 980 5132
rect 1044 5130 1050 5132
rect 5165 5130 5231 5133
rect 9622 5130 9628 5132
rect 1044 5128 5231 5130
rect 1044 5072 5170 5128
rect 5226 5072 5231 5128
rect 1044 5070 5231 5072
rect 1044 5068 1050 5070
rect 5165 5067 5231 5070
rect 5398 5070 9628 5130
rect 3969 4994 4035 4997
rect 5398 4994 5458 5070
rect 9622 5068 9628 5070
rect 9692 5068 9698 5132
rect 11010 5130 11070 5206
rect 11513 5264 13308 5266
rect 11513 5208 11518 5264
rect 11574 5208 13308 5264
rect 11513 5206 13308 5208
rect 11513 5203 11579 5206
rect 13302 5204 13308 5206
rect 13372 5204 13378 5268
rect 14549 5130 14615 5133
rect 11010 5128 14615 5130
rect 11010 5072 14554 5128
rect 14610 5072 14615 5128
rect 11010 5070 14615 5072
rect 14549 5067 14615 5070
rect 3969 4992 5458 4994
rect 3969 4936 3974 4992
rect 4030 4936 5458 4992
rect 3969 4934 5458 4936
rect 3969 4931 4035 4934
rect 6310 4932 6316 4996
rect 6380 4994 6386 4996
rect 6729 4994 6795 4997
rect 6380 4992 6795 4994
rect 6380 4936 6734 4992
rect 6790 4936 6795 4992
rect 6380 4934 6795 4936
rect 6380 4932 6386 4934
rect 6729 4931 6795 4934
rect 7414 4932 7420 4996
rect 7484 4994 7490 4996
rect 10777 4994 10843 4997
rect 7484 4992 10843 4994
rect 7484 4936 10782 4992
rect 10838 4936 10843 4992
rect 7484 4934 10843 4936
rect 7484 4932 7490 4934
rect 10777 4931 10843 4934
rect 1946 4928 2262 4929
rect 1946 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2262 4928
rect 1946 4863 2262 4864
rect 6946 4928 7262 4929
rect 6946 4864 6952 4928
rect 7016 4864 7032 4928
rect 7096 4864 7112 4928
rect 7176 4864 7192 4928
rect 7256 4864 7262 4928
rect 6946 4863 7262 4864
rect 11946 4928 12262 4929
rect 11946 4864 11952 4928
rect 12016 4864 12032 4928
rect 12096 4864 12112 4928
rect 12176 4864 12192 4928
rect 12256 4864 12262 4928
rect 11946 4863 12262 4864
rect 16946 4928 17262 4929
rect 16946 4864 16952 4928
rect 17016 4864 17032 4928
rect 17096 4864 17112 4928
rect 17176 4864 17192 4928
rect 17256 4864 17262 4928
rect 16946 4863 17262 4864
rect 2773 4858 2839 4861
rect 5206 4858 5212 4860
rect 2773 4856 5212 4858
rect 2773 4800 2778 4856
rect 2834 4800 5212 4856
rect 2773 4798 5212 4800
rect 2773 4795 2839 4798
rect 5206 4796 5212 4798
rect 5276 4796 5282 4860
rect 12433 4858 12499 4861
rect 13629 4858 13695 4861
rect 14825 4860 14891 4861
rect 12433 4856 13695 4858
rect 12433 4800 12438 4856
rect 12494 4800 13634 4856
rect 13690 4800 13695 4856
rect 12433 4798 13695 4800
rect 12433 4795 12499 4798
rect 13629 4795 13695 4798
rect 14774 4796 14780 4860
rect 14844 4858 14891 4860
rect 14844 4856 14936 4858
rect 14886 4800 14936 4856
rect 14844 4798 14936 4800
rect 14844 4796 14891 4798
rect 14825 4795 14891 4796
rect 4797 4722 4863 4725
rect 6637 4722 6703 4725
rect 14641 4722 14707 4725
rect 15142 4722 15148 4724
rect 4797 4720 14520 4722
rect 4797 4664 4802 4720
rect 4858 4664 6642 4720
rect 6698 4664 14520 4720
rect 4797 4662 14520 4664
rect 4797 4659 4863 4662
rect 6637 4659 6703 4662
rect 4705 4586 4771 4589
rect 5022 4586 5028 4588
rect 4705 4584 5028 4586
rect 4705 4528 4710 4584
rect 4766 4528 5028 4584
rect 4705 4526 5028 4528
rect 4705 4523 4771 4526
rect 5022 4524 5028 4526
rect 5092 4524 5098 4588
rect 5441 4586 5507 4589
rect 7925 4586 7991 4589
rect 9673 4586 9739 4589
rect 5441 4584 7991 4586
rect 5441 4528 5446 4584
rect 5502 4528 7930 4584
rect 7986 4528 7991 4584
rect 5441 4526 7991 4528
rect 5441 4523 5507 4526
rect 7925 4523 7991 4526
rect 8388 4584 9739 4586
rect 8388 4528 9678 4584
rect 9734 4528 9739 4584
rect 8388 4526 9739 4528
rect 8388 4453 8448 4526
rect 9673 4523 9739 4526
rect 11789 4586 11855 4589
rect 12985 4586 13051 4589
rect 11789 4584 13051 4586
rect 11789 4528 11794 4584
rect 11850 4528 12990 4584
rect 13046 4528 13051 4584
rect 11789 4526 13051 4528
rect 14460 4586 14520 4662
rect 14641 4720 15148 4722
rect 14641 4664 14646 4720
rect 14702 4664 15148 4720
rect 14641 4662 15148 4664
rect 14641 4659 14707 4662
rect 15142 4660 15148 4662
rect 15212 4660 15218 4724
rect 16430 4586 16436 4588
rect 14460 4526 16436 4586
rect 11789 4523 11855 4526
rect 12985 4523 13051 4526
rect 16254 4453 16314 4526
rect 16430 4524 16436 4526
rect 16500 4524 16506 4588
rect 5809 4450 5875 4453
rect 6126 4450 6132 4452
rect 5809 4448 6132 4450
rect 5809 4392 5814 4448
rect 5870 4392 6132 4448
rect 5809 4390 6132 4392
rect 5809 4387 5875 4390
rect 6126 4388 6132 4390
rect 6196 4388 6202 4452
rect 6637 4450 6703 4453
rect 7414 4450 7420 4452
rect 6637 4448 7420 4450
rect 6637 4392 6642 4448
rect 6698 4392 7420 4448
rect 6637 4390 7420 4392
rect 6637 4387 6703 4390
rect 7414 4388 7420 4390
rect 7484 4388 7490 4452
rect 8385 4448 8451 4453
rect 8385 4392 8390 4448
rect 8446 4392 8451 4448
rect 8385 4387 8451 4392
rect 8845 4450 8911 4453
rect 12433 4450 12499 4453
rect 13537 4452 13603 4453
rect 13486 4450 13492 4452
rect 8845 4448 12499 4450
rect 8845 4392 8850 4448
rect 8906 4392 12438 4448
rect 12494 4392 12499 4448
rect 8845 4390 12499 4392
rect 13446 4390 13492 4450
rect 13556 4448 13603 4452
rect 13598 4392 13603 4448
rect 8845 4387 8911 4390
rect 12433 4387 12499 4390
rect 13486 4388 13492 4390
rect 13556 4388 13603 4392
rect 13670 4388 13676 4452
rect 13740 4450 13746 4452
rect 15929 4450 15995 4453
rect 13740 4448 15995 4450
rect 13740 4392 15934 4448
rect 15990 4392 15995 4448
rect 13740 4390 15995 4392
rect 16254 4448 16363 4453
rect 16254 4392 16302 4448
rect 16358 4392 16363 4448
rect 16254 4390 16363 4392
rect 13740 4388 13746 4390
rect 13537 4387 13603 4388
rect 15929 4387 15995 4390
rect 16297 4387 16363 4390
rect 2606 4384 2922 4385
rect 2606 4320 2612 4384
rect 2676 4320 2692 4384
rect 2756 4320 2772 4384
rect 2836 4320 2852 4384
rect 2916 4320 2922 4384
rect 2606 4319 2922 4320
rect 7606 4384 7922 4385
rect 7606 4320 7612 4384
rect 7676 4320 7692 4384
rect 7756 4320 7772 4384
rect 7836 4320 7852 4384
rect 7916 4320 7922 4384
rect 7606 4319 7922 4320
rect 12606 4384 12922 4385
rect 12606 4320 12612 4384
rect 12676 4320 12692 4384
rect 12756 4320 12772 4384
rect 12836 4320 12852 4384
rect 12916 4320 12922 4384
rect 12606 4319 12922 4320
rect 17606 4384 17922 4385
rect 17606 4320 17612 4384
rect 17676 4320 17692 4384
rect 17756 4320 17772 4384
rect 17836 4320 17852 4384
rect 17916 4320 17922 4384
rect 17606 4319 17922 4320
rect 3182 4252 3188 4316
rect 3252 4314 3258 4316
rect 3325 4314 3391 4317
rect 6085 4314 6151 4317
rect 7373 4314 7439 4317
rect 11094 4314 11100 4316
rect 3252 4312 6010 4314
rect 3252 4256 3330 4312
rect 3386 4256 6010 4312
rect 3252 4254 6010 4256
rect 3252 4252 3258 4254
rect 3325 4251 3391 4254
rect 1393 4178 1459 4181
rect 5441 4178 5507 4181
rect 1393 4176 5507 4178
rect 1393 4120 1398 4176
rect 1454 4120 5446 4176
rect 5502 4120 5507 4176
rect 1393 4118 5507 4120
rect 5950 4178 6010 4254
rect 6085 4312 7439 4314
rect 6085 4256 6090 4312
rect 6146 4256 7378 4312
rect 7434 4256 7439 4312
rect 6085 4254 7439 4256
rect 6085 4251 6151 4254
rect 7373 4251 7439 4254
rect 9446 4254 11100 4314
rect 7189 4178 7255 4181
rect 8334 4178 8340 4180
rect 5950 4176 8340 4178
rect 5950 4120 7194 4176
rect 7250 4120 8340 4176
rect 5950 4118 8340 4120
rect 1393 4115 1459 4118
rect 5441 4115 5507 4118
rect 7189 4115 7255 4118
rect 8334 4116 8340 4118
rect 8404 4116 8410 4180
rect 1209 4042 1275 4045
rect 3877 4042 3943 4045
rect 1209 4040 3943 4042
rect 1209 3984 1214 4040
rect 1270 3984 3882 4040
rect 3938 3984 3943 4040
rect 1209 3982 3943 3984
rect 1209 3979 1275 3982
rect 3877 3979 3943 3982
rect 4981 4042 5047 4045
rect 8385 4042 8451 4045
rect 4981 4040 8451 4042
rect 4981 3984 4986 4040
rect 5042 3984 8390 4040
rect 8446 3984 8451 4040
rect 4981 3982 8451 3984
rect 4981 3979 5047 3982
rect 8385 3979 8451 3982
rect 8845 4042 8911 4045
rect 9446 4042 9506 4254
rect 11094 4252 11100 4254
rect 11164 4252 11170 4316
rect 9673 4178 9739 4181
rect 12341 4178 12407 4181
rect 14958 4178 14964 4180
rect 9673 4176 12082 4178
rect 9673 4120 9678 4176
rect 9734 4120 12082 4176
rect 9673 4118 12082 4120
rect 9673 4115 9739 4118
rect 8845 4040 9506 4042
rect 8845 3984 8850 4040
rect 8906 3984 9506 4040
rect 8845 3982 9506 3984
rect 9581 4042 9647 4045
rect 10726 4042 10732 4044
rect 9581 4040 10732 4042
rect 9581 3984 9586 4040
rect 9642 3984 10732 4040
rect 9581 3982 10732 3984
rect 8845 3979 8911 3982
rect 9581 3979 9647 3982
rect 10726 3980 10732 3982
rect 10796 3980 10802 4044
rect 10961 4042 11027 4045
rect 11646 4042 11652 4044
rect 10961 4040 11652 4042
rect 10961 3984 10966 4040
rect 11022 3984 11652 4040
rect 10961 3982 11652 3984
rect 10961 3979 11027 3982
rect 11646 3980 11652 3982
rect 11716 3980 11722 4044
rect 12022 4042 12082 4118
rect 12341 4176 14964 4178
rect 12341 4120 12346 4176
rect 12402 4120 14964 4176
rect 12341 4118 14964 4120
rect 12341 4115 12407 4118
rect 14958 4116 14964 4118
rect 15028 4116 15034 4180
rect 15142 4116 15148 4180
rect 15212 4178 15218 4180
rect 15653 4178 15719 4181
rect 15212 4176 15719 4178
rect 15212 4120 15658 4176
rect 15714 4120 15719 4176
rect 15212 4118 15719 4120
rect 15212 4116 15218 4118
rect 15653 4115 15719 4118
rect 16021 4180 16087 4181
rect 16021 4176 16068 4180
rect 16132 4178 16138 4180
rect 16021 4120 16026 4176
rect 16021 4116 16068 4120
rect 16132 4118 16178 4178
rect 16132 4116 16138 4118
rect 16021 4115 16087 4116
rect 14038 4042 14044 4044
rect 12022 3982 14044 4042
rect 14038 3980 14044 3982
rect 14108 3980 14114 4044
rect 18229 4042 18295 4045
rect 18822 4042 18828 4044
rect 18229 4040 18828 4042
rect 18229 3984 18234 4040
rect 18290 3984 18828 4040
rect 18229 3982 18828 3984
rect 18229 3979 18295 3982
rect 18822 3980 18828 3982
rect 18892 3980 18898 4044
rect 0 3906 800 3936
rect 1393 3906 1459 3909
rect 0 3904 1459 3906
rect 0 3848 1398 3904
rect 1454 3848 1459 3904
rect 0 3846 1459 3848
rect 0 3816 800 3846
rect 1393 3843 1459 3846
rect 2405 3906 2471 3909
rect 4337 3906 4403 3909
rect 2405 3904 4403 3906
rect 2405 3848 2410 3904
rect 2466 3848 4342 3904
rect 4398 3848 4403 3904
rect 2405 3846 4403 3848
rect 2405 3843 2471 3846
rect 4337 3843 4403 3846
rect 4470 3844 4476 3908
rect 4540 3906 4546 3908
rect 4981 3906 5047 3909
rect 4540 3904 5047 3906
rect 4540 3848 4986 3904
rect 5042 3848 5047 3904
rect 4540 3846 5047 3848
rect 4540 3844 4546 3846
rect 4981 3843 5047 3846
rect 5901 3906 5967 3909
rect 8569 3908 8635 3909
rect 6310 3906 6316 3908
rect 5901 3904 6316 3906
rect 5901 3848 5906 3904
rect 5962 3848 6316 3904
rect 5901 3846 6316 3848
rect 5901 3843 5967 3846
rect 6310 3844 6316 3846
rect 6380 3844 6386 3908
rect 8518 3844 8524 3908
rect 8588 3906 8635 3908
rect 8937 3906 9003 3909
rect 11697 3906 11763 3909
rect 8588 3904 8680 3906
rect 8630 3848 8680 3904
rect 8588 3846 8680 3848
rect 8937 3904 11763 3906
rect 8937 3848 8942 3904
rect 8998 3848 11702 3904
rect 11758 3848 11763 3904
rect 8937 3846 11763 3848
rect 8588 3844 8635 3846
rect 8569 3843 8635 3844
rect 8937 3843 9003 3846
rect 11697 3843 11763 3846
rect 18413 3906 18479 3909
rect 19200 3906 20000 3936
rect 18413 3904 20000 3906
rect 18413 3848 18418 3904
rect 18474 3848 20000 3904
rect 18413 3846 20000 3848
rect 18413 3843 18479 3846
rect 1946 3840 2262 3841
rect 1946 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2262 3840
rect 1946 3775 2262 3776
rect 6946 3840 7262 3841
rect 6946 3776 6952 3840
rect 7016 3776 7032 3840
rect 7096 3776 7112 3840
rect 7176 3776 7192 3840
rect 7256 3776 7262 3840
rect 6946 3775 7262 3776
rect 11946 3840 12262 3841
rect 11946 3776 11952 3840
rect 12016 3776 12032 3840
rect 12096 3776 12112 3840
rect 12176 3776 12192 3840
rect 12256 3776 12262 3840
rect 11946 3775 12262 3776
rect 16946 3840 17262 3841
rect 16946 3776 16952 3840
rect 17016 3776 17032 3840
rect 17096 3776 17112 3840
rect 17176 3776 17192 3840
rect 17256 3776 17262 3840
rect 19200 3816 20000 3846
rect 16946 3775 17262 3776
rect 4613 3770 4679 3773
rect 6453 3770 6519 3773
rect 9254 3770 9260 3772
rect 4613 3768 6519 3770
rect 4613 3712 4618 3768
rect 4674 3712 6458 3768
rect 6514 3712 6519 3768
rect 4613 3710 6519 3712
rect 4613 3707 4679 3710
rect 6453 3707 6519 3710
rect 7376 3710 9260 3770
rect 933 3634 999 3637
rect 5441 3634 5507 3637
rect 5942 3634 5948 3636
rect 933 3632 4722 3634
rect 933 3576 938 3632
rect 994 3576 4722 3632
rect 933 3574 4722 3576
rect 933 3571 999 3574
rect 3049 3498 3115 3501
rect 3366 3498 3372 3500
rect 3049 3496 3372 3498
rect 3049 3440 3054 3496
rect 3110 3440 3372 3496
rect 3049 3438 3372 3440
rect 3049 3435 3115 3438
rect 3366 3436 3372 3438
rect 3436 3436 3442 3500
rect 4102 3436 4108 3500
rect 4172 3498 4178 3500
rect 4521 3498 4587 3501
rect 4172 3496 4587 3498
rect 4172 3440 4526 3496
rect 4582 3440 4587 3496
rect 4172 3438 4587 3440
rect 4662 3498 4722 3574
rect 5441 3632 5948 3634
rect 5441 3576 5446 3632
rect 5502 3576 5948 3632
rect 5441 3574 5948 3576
rect 5441 3571 5507 3574
rect 5942 3572 5948 3574
rect 6012 3634 6018 3636
rect 7005 3634 7071 3637
rect 6012 3632 7071 3634
rect 6012 3576 7010 3632
rect 7066 3576 7071 3632
rect 6012 3574 7071 3576
rect 6012 3572 6018 3574
rect 7005 3571 7071 3574
rect 7189 3634 7255 3637
rect 7376 3634 7436 3710
rect 9254 3708 9260 3710
rect 9324 3708 9330 3772
rect 12341 3770 12407 3773
rect 12341 3768 16268 3770
rect 12341 3712 12346 3768
rect 12402 3712 16268 3768
rect 12341 3710 16268 3712
rect 12341 3707 12407 3710
rect 7189 3632 7436 3634
rect 7189 3576 7194 3632
rect 7250 3576 7436 3632
rect 7189 3574 7436 3576
rect 8201 3634 8267 3637
rect 11697 3634 11763 3637
rect 8201 3632 11763 3634
rect 8201 3576 8206 3632
rect 8262 3576 11702 3632
rect 11758 3576 11763 3632
rect 8201 3574 11763 3576
rect 7189 3571 7255 3574
rect 8201 3571 8267 3574
rect 11697 3571 11763 3574
rect 12801 3634 12867 3637
rect 13854 3634 13860 3636
rect 12801 3632 13860 3634
rect 12801 3576 12806 3632
rect 12862 3576 13860 3632
rect 12801 3574 13860 3576
rect 12801 3571 12867 3574
rect 13854 3572 13860 3574
rect 13924 3572 13930 3636
rect 16208 3634 16268 3710
rect 17953 3634 18019 3637
rect 16208 3632 18019 3634
rect 16208 3576 17958 3632
rect 18014 3576 18019 3632
rect 16208 3574 18019 3576
rect 17953 3571 18019 3574
rect 5625 3498 5691 3501
rect 4662 3496 5691 3498
rect 4662 3440 5630 3496
rect 5686 3440 5691 3496
rect 4662 3438 5691 3440
rect 4172 3436 4178 3438
rect 4521 3435 4587 3438
rect 5625 3435 5691 3438
rect 6085 3498 6151 3501
rect 18137 3498 18203 3501
rect 6085 3496 18203 3498
rect 6085 3440 6090 3496
rect 6146 3440 18142 3496
rect 18198 3440 18203 3496
rect 6085 3438 18203 3440
rect 6085 3435 6151 3438
rect 18137 3435 18203 3438
rect 3417 3362 3483 3365
rect 5533 3362 5599 3365
rect 3417 3360 5599 3362
rect 3417 3304 3422 3360
rect 3478 3304 5538 3360
rect 5594 3304 5599 3360
rect 3417 3302 5599 3304
rect 3417 3299 3483 3302
rect 5533 3299 5599 3302
rect 6494 3300 6500 3364
rect 6564 3362 6570 3364
rect 7281 3362 7347 3365
rect 6564 3360 7347 3362
rect 6564 3304 7286 3360
rect 7342 3304 7347 3360
rect 6564 3302 7347 3304
rect 6564 3300 6570 3302
rect 7281 3299 7347 3302
rect 9254 3300 9260 3364
rect 9324 3362 9330 3364
rect 12341 3362 12407 3365
rect 9324 3360 12407 3362
rect 9324 3304 12346 3360
rect 12402 3304 12407 3360
rect 9324 3302 12407 3304
rect 9324 3300 9330 3302
rect 12341 3299 12407 3302
rect 16113 3362 16179 3365
rect 16573 3362 16639 3365
rect 16849 3364 16915 3365
rect 16798 3362 16804 3364
rect 16113 3360 16639 3362
rect 16113 3304 16118 3360
rect 16174 3304 16578 3360
rect 16634 3304 16639 3360
rect 16113 3302 16639 3304
rect 16758 3302 16804 3362
rect 16868 3360 16915 3364
rect 16910 3304 16915 3360
rect 16113 3299 16179 3302
rect 16573 3299 16639 3302
rect 16798 3300 16804 3302
rect 16868 3300 16915 3304
rect 16849 3299 16915 3300
rect 2606 3296 2922 3297
rect 2606 3232 2612 3296
rect 2676 3232 2692 3296
rect 2756 3232 2772 3296
rect 2836 3232 2852 3296
rect 2916 3232 2922 3296
rect 2606 3231 2922 3232
rect 7606 3296 7922 3297
rect 7606 3232 7612 3296
rect 7676 3232 7692 3296
rect 7756 3232 7772 3296
rect 7836 3232 7852 3296
rect 7916 3232 7922 3296
rect 7606 3231 7922 3232
rect 12606 3296 12922 3297
rect 12606 3232 12612 3296
rect 12676 3232 12692 3296
rect 12756 3232 12772 3296
rect 12836 3232 12852 3296
rect 12916 3232 12922 3296
rect 12606 3231 12922 3232
rect 17606 3296 17922 3297
rect 17606 3232 17612 3296
rect 17676 3232 17692 3296
rect 17756 3232 17772 3296
rect 17836 3232 17852 3296
rect 17916 3232 17922 3296
rect 17606 3231 17922 3232
rect 8293 3226 8359 3229
rect 9489 3226 9555 3229
rect 8293 3224 9555 3226
rect 8293 3168 8298 3224
rect 8354 3168 9494 3224
rect 9550 3168 9555 3224
rect 8293 3166 9555 3168
rect 8293 3163 8359 3166
rect 9489 3163 9555 3166
rect 11278 3164 11284 3228
rect 11348 3226 11354 3228
rect 12433 3226 12499 3229
rect 11348 3224 12499 3226
rect 11348 3168 12438 3224
rect 12494 3168 12499 3224
rect 11348 3166 12499 3168
rect 11348 3164 11354 3166
rect 12433 3163 12499 3166
rect 2773 3090 2839 3093
rect 3734 3090 3740 3092
rect 2773 3088 3740 3090
rect 2773 3032 2778 3088
rect 2834 3032 3740 3088
rect 2773 3030 3740 3032
rect 2773 3027 2839 3030
rect 3734 3028 3740 3030
rect 3804 3028 3810 3092
rect 4981 3090 5047 3093
rect 15377 3090 15443 3093
rect 4981 3088 15443 3090
rect 4981 3032 4986 3088
rect 5042 3032 15382 3088
rect 15438 3032 15443 3088
rect 4981 3030 15443 3032
rect 4981 3027 5047 3030
rect 15377 3027 15443 3030
rect 2446 2892 2452 2956
rect 2516 2954 2522 2956
rect 7925 2954 7991 2957
rect 2516 2952 7991 2954
rect 2516 2896 7930 2952
rect 7986 2896 7991 2952
rect 2516 2894 7991 2896
rect 2516 2892 2522 2894
rect 7925 2891 7991 2894
rect 8293 2954 8359 2957
rect 9857 2954 9923 2957
rect 8293 2952 9923 2954
rect 8293 2896 8298 2952
rect 8354 2896 9862 2952
rect 9918 2896 9923 2952
rect 8293 2894 9923 2896
rect 8293 2891 8359 2894
rect 9857 2891 9923 2894
rect 10777 2954 10843 2957
rect 15561 2954 15627 2957
rect 10777 2952 15627 2954
rect 10777 2896 10782 2952
rect 10838 2896 15566 2952
rect 15622 2896 15627 2952
rect 10777 2894 15627 2896
rect 10777 2891 10843 2894
rect 15561 2891 15627 2894
rect 8845 2818 8911 2821
rect 7652 2816 8911 2818
rect 7652 2760 8850 2816
rect 8906 2760 8911 2816
rect 7652 2758 8911 2760
rect 1946 2752 2262 2753
rect 1946 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2262 2752
rect 1946 2687 2262 2688
rect 6946 2752 7262 2753
rect 6946 2688 6952 2752
rect 7016 2688 7032 2752
rect 7096 2688 7112 2752
rect 7176 2688 7192 2752
rect 7256 2688 7262 2752
rect 6946 2687 7262 2688
rect 3550 2620 3556 2684
rect 3620 2682 3626 2684
rect 6545 2682 6611 2685
rect 3620 2680 6611 2682
rect 3620 2624 6550 2680
rect 6606 2624 6611 2680
rect 3620 2622 6611 2624
rect 3620 2620 3626 2622
rect 6545 2619 6611 2622
rect 1342 2484 1348 2548
rect 1412 2546 1418 2548
rect 7652 2546 7712 2758
rect 8845 2755 8911 2758
rect 11946 2752 12262 2753
rect 11946 2688 11952 2752
rect 12016 2688 12032 2752
rect 12096 2688 12112 2752
rect 12176 2688 12192 2752
rect 12256 2688 12262 2752
rect 11946 2687 12262 2688
rect 16946 2752 17262 2753
rect 16946 2688 16952 2752
rect 17016 2688 17032 2752
rect 17096 2688 17112 2752
rect 17176 2688 17192 2752
rect 17256 2688 17262 2752
rect 16946 2687 17262 2688
rect 8201 2684 8267 2685
rect 8150 2682 8156 2684
rect 8110 2622 8156 2682
rect 8220 2680 8267 2684
rect 8262 2624 8267 2680
rect 8150 2620 8156 2622
rect 8220 2620 8267 2624
rect 8201 2619 8267 2620
rect 8661 2684 8727 2685
rect 8661 2680 8708 2684
rect 8772 2682 8778 2684
rect 8661 2624 8666 2680
rect 8661 2620 8708 2624
rect 8772 2622 8818 2682
rect 8772 2620 8778 2622
rect 8886 2620 8892 2684
rect 8956 2682 8962 2684
rect 9029 2682 9095 2685
rect 8956 2680 9095 2682
rect 8956 2624 9034 2680
rect 9090 2624 9095 2680
rect 8956 2622 9095 2624
rect 8956 2620 8962 2622
rect 8661 2619 8727 2620
rect 9029 2619 9095 2622
rect 13721 2682 13787 2685
rect 16246 2682 16252 2684
rect 13721 2680 16252 2682
rect 13721 2624 13726 2680
rect 13782 2624 16252 2680
rect 13721 2622 16252 2624
rect 13721 2619 13787 2622
rect 16246 2620 16252 2622
rect 16316 2620 16322 2684
rect 1412 2486 7712 2546
rect 8569 2546 8635 2549
rect 10358 2546 10364 2548
rect 8569 2544 10364 2546
rect 8569 2488 8574 2544
rect 8630 2488 10364 2544
rect 8569 2486 10364 2488
rect 1412 2484 1418 2486
rect 8569 2483 8635 2486
rect 10358 2484 10364 2486
rect 10428 2484 10434 2548
rect 10910 2484 10916 2548
rect 10980 2546 10986 2548
rect 11973 2546 12039 2549
rect 10980 2544 12039 2546
rect 10980 2488 11978 2544
rect 12034 2488 12039 2544
rect 10980 2486 12039 2488
rect 10980 2484 10986 2486
rect 11973 2483 12039 2486
rect 16614 2484 16620 2548
rect 16684 2546 16690 2548
rect 16941 2546 17007 2549
rect 16684 2544 17007 2546
rect 16684 2488 16946 2544
rect 17002 2488 17007 2544
rect 16684 2486 17007 2488
rect 16684 2484 16690 2486
rect 16941 2483 17007 2486
rect 1485 2410 1551 2413
rect 8477 2410 8543 2413
rect 1485 2408 8543 2410
rect 1485 2352 1490 2408
rect 1546 2352 8482 2408
rect 8538 2352 8543 2408
rect 1485 2350 8543 2352
rect 1485 2347 1551 2350
rect 8477 2347 8543 2350
rect 11329 2410 11395 2413
rect 14406 2410 14412 2412
rect 11329 2408 14412 2410
rect 11329 2352 11334 2408
rect 11390 2352 14412 2408
rect 11329 2350 14412 2352
rect 11329 2347 11395 2350
rect 14406 2348 14412 2350
rect 14476 2348 14482 2412
rect 17953 2410 18019 2413
rect 18638 2410 18644 2412
rect 17953 2408 18644 2410
rect 17953 2352 17958 2408
rect 18014 2352 18644 2408
rect 17953 2350 18644 2352
rect 17953 2347 18019 2350
rect 18638 2348 18644 2350
rect 18708 2348 18714 2412
rect 5390 2212 5396 2276
rect 5460 2274 5466 2276
rect 7465 2274 7531 2277
rect 5460 2272 7531 2274
rect 5460 2216 7470 2272
rect 7526 2216 7531 2272
rect 5460 2214 7531 2216
rect 5460 2212 5466 2214
rect 7465 2211 7531 2214
rect 8017 2274 8083 2277
rect 8017 2272 12450 2274
rect 8017 2216 8022 2272
rect 8078 2216 12450 2272
rect 8017 2214 12450 2216
rect 8017 2211 8083 2214
rect 2606 2208 2922 2209
rect 2606 2144 2612 2208
rect 2676 2144 2692 2208
rect 2756 2144 2772 2208
rect 2836 2144 2852 2208
rect 2916 2144 2922 2208
rect 2606 2143 2922 2144
rect 7606 2208 7922 2209
rect 7606 2144 7612 2208
rect 7676 2144 7692 2208
rect 7756 2144 7772 2208
rect 7836 2144 7852 2208
rect 7916 2144 7922 2208
rect 7606 2143 7922 2144
rect 3233 2138 3299 2141
rect 3233 2136 5826 2138
rect 3233 2080 3238 2136
rect 3294 2080 5826 2136
rect 3233 2078 5826 2080
rect 3233 2075 3299 2078
rect 5766 2002 5826 2078
rect 12390 2002 12450 2214
rect 12606 2208 12922 2209
rect 12606 2144 12612 2208
rect 12676 2144 12692 2208
rect 12756 2144 12772 2208
rect 12836 2144 12852 2208
rect 12916 2144 12922 2208
rect 12606 2143 12922 2144
rect 17606 2208 17922 2209
rect 17606 2144 17612 2208
rect 17676 2144 17692 2208
rect 17756 2144 17772 2208
rect 17836 2144 17852 2208
rect 17916 2144 17922 2208
rect 17606 2143 17922 2144
rect 15326 2002 15332 2004
rect 5766 1942 10794 2002
rect 12390 1942 15332 2002
rect 6085 1866 6151 1869
rect 10542 1866 10548 1868
rect 6085 1864 10548 1866
rect 6085 1808 6090 1864
rect 6146 1808 10548 1864
rect 6085 1806 10548 1808
rect 6085 1803 6151 1806
rect 10542 1804 10548 1806
rect 10612 1804 10618 1868
rect 10734 1866 10794 1942
rect 15326 1940 15332 1942
rect 15396 1940 15402 2004
rect 10734 1806 12450 1866
rect 10317 1730 10383 1733
rect 2730 1728 10383 1730
rect 2730 1672 10322 1728
rect 10378 1672 10383 1728
rect 2730 1670 10383 1672
rect 12390 1730 12450 1806
rect 16665 1730 16731 1733
rect 12390 1728 16731 1730
rect 12390 1672 16670 1728
rect 16726 1672 16731 1728
rect 12390 1670 16731 1672
rect 0 1458 800 1488
rect 2405 1458 2471 1461
rect 0 1456 2471 1458
rect 0 1400 2410 1456
rect 2466 1400 2471 1456
rect 0 1398 2471 1400
rect 0 1368 800 1398
rect 2405 1395 2471 1398
rect 2589 1458 2655 1461
rect 2730 1458 2790 1670
rect 10317 1667 10383 1670
rect 16665 1667 16731 1670
rect 17902 1668 17908 1732
rect 17972 1730 17978 1732
rect 19006 1730 19012 1732
rect 17972 1670 19012 1730
rect 17972 1668 17978 1670
rect 19006 1668 19012 1670
rect 19076 1668 19082 1732
rect 6545 1594 6611 1597
rect 18229 1594 18295 1597
rect 6545 1592 18295 1594
rect 6545 1536 6550 1592
rect 6606 1536 18234 1592
rect 18290 1536 18295 1592
rect 6545 1534 18295 1536
rect 6545 1531 6611 1534
rect 18229 1531 18295 1534
rect 2589 1456 2790 1458
rect 2589 1400 2594 1456
rect 2650 1400 2790 1456
rect 2589 1398 2790 1400
rect 7189 1458 7255 1461
rect 17902 1458 17908 1460
rect 7189 1456 17908 1458
rect 7189 1400 7194 1456
rect 7250 1400 17908 1456
rect 7189 1398 17908 1400
rect 2589 1395 2655 1398
rect 7189 1395 7255 1398
rect 17902 1396 17908 1398
rect 17972 1396 17978 1460
rect 18321 1458 18387 1461
rect 19200 1458 20000 1488
rect 18321 1456 20000 1458
rect 18321 1400 18326 1456
rect 18382 1400 20000 1456
rect 18321 1398 20000 1400
rect 18321 1395 18387 1398
rect 19200 1368 20000 1398
rect 4797 1186 4863 1189
rect 8385 1186 8451 1189
rect 4797 1184 8451 1186
rect 4797 1128 4802 1184
rect 4858 1128 8390 1184
rect 8446 1128 8451 1184
rect 4797 1126 8451 1128
rect 4797 1123 4863 1126
rect 8385 1123 8451 1126
rect 1393 1050 1459 1053
rect 1710 1050 1716 1052
rect 1393 1048 1716 1050
rect 1393 992 1398 1048
rect 1454 992 1716 1048
rect 1393 990 1716 992
rect 1393 987 1459 990
rect 1710 988 1716 990
rect 1780 988 1786 1052
rect 7373 1050 7439 1053
rect 15285 1050 15351 1053
rect 7373 1048 15351 1050
rect 7373 992 7378 1048
rect 7434 992 15290 1048
rect 15346 992 15351 1048
rect 7373 990 15351 992
rect 7373 987 7439 990
rect 15285 987 15351 990
rect 3918 852 3924 916
rect 3988 914 3994 916
rect 15837 914 15903 917
rect 3988 912 15903 914
rect 3988 856 15842 912
rect 15898 856 15903 912
rect 3988 854 15903 856
rect 3988 852 3994 854
rect 15837 851 15903 854
rect 790 716 796 780
rect 860 778 866 780
rect 12341 778 12407 781
rect 860 776 12407 778
rect 860 720 12346 776
rect 12402 720 12407 776
rect 860 718 12407 720
rect 860 716 866 718
rect 12341 715 12407 718
rect 4654 580 4660 644
rect 4724 642 4730 644
rect 11605 642 11671 645
rect 4724 640 11671 642
rect 4724 584 11610 640
rect 11666 584 11671 640
rect 4724 582 11671 584
rect 4724 580 4730 582
rect 11605 579 11671 582
rect 3877 506 3943 509
rect 13118 506 13124 508
rect 3877 504 13124 506
rect 3877 448 3882 504
rect 3938 448 13124 504
rect 3877 446 13124 448
rect 3877 443 3943 446
rect 13118 444 13124 446
rect 13188 444 13194 508
<< via3 >>
rect 15884 18668 15948 18732
rect 5028 18532 5092 18596
rect 1532 18396 1596 18460
rect 13860 18260 13924 18324
rect 14596 18124 14660 18188
rect 5764 18048 5828 18052
rect 5764 17992 5814 18048
rect 5814 17992 5828 18048
rect 5764 17988 5828 17992
rect 13492 17580 13556 17644
rect 2612 17436 2676 17440
rect 2612 17380 2616 17436
rect 2616 17380 2672 17436
rect 2672 17380 2676 17436
rect 2612 17376 2676 17380
rect 2692 17436 2756 17440
rect 2692 17380 2696 17436
rect 2696 17380 2752 17436
rect 2752 17380 2756 17436
rect 2692 17376 2756 17380
rect 2772 17436 2836 17440
rect 2772 17380 2776 17436
rect 2776 17380 2832 17436
rect 2832 17380 2836 17436
rect 2772 17376 2836 17380
rect 2852 17436 2916 17440
rect 2852 17380 2856 17436
rect 2856 17380 2912 17436
rect 2912 17380 2916 17436
rect 2852 17376 2916 17380
rect 7612 17436 7676 17440
rect 7612 17380 7616 17436
rect 7616 17380 7672 17436
rect 7672 17380 7676 17436
rect 7612 17376 7676 17380
rect 7692 17436 7756 17440
rect 7692 17380 7696 17436
rect 7696 17380 7752 17436
rect 7752 17380 7756 17436
rect 7692 17376 7756 17380
rect 7772 17436 7836 17440
rect 7772 17380 7776 17436
rect 7776 17380 7832 17436
rect 7832 17380 7836 17436
rect 7772 17376 7836 17380
rect 7852 17436 7916 17440
rect 7852 17380 7856 17436
rect 7856 17380 7912 17436
rect 7912 17380 7916 17436
rect 7852 17376 7916 17380
rect 12612 17436 12676 17440
rect 12612 17380 12616 17436
rect 12616 17380 12672 17436
rect 12672 17380 12676 17436
rect 12612 17376 12676 17380
rect 12692 17436 12756 17440
rect 12692 17380 12696 17436
rect 12696 17380 12752 17436
rect 12752 17380 12756 17436
rect 12692 17376 12756 17380
rect 12772 17436 12836 17440
rect 12772 17380 12776 17436
rect 12776 17380 12832 17436
rect 12832 17380 12836 17436
rect 12772 17376 12836 17380
rect 12852 17436 12916 17440
rect 12852 17380 12856 17436
rect 12856 17380 12912 17436
rect 12912 17380 12916 17436
rect 12852 17376 12916 17380
rect 17612 17436 17676 17440
rect 17612 17380 17616 17436
rect 17616 17380 17672 17436
rect 17672 17380 17676 17436
rect 17612 17376 17676 17380
rect 17692 17436 17756 17440
rect 17692 17380 17696 17436
rect 17696 17380 17752 17436
rect 17752 17380 17756 17436
rect 17692 17376 17756 17380
rect 17772 17436 17836 17440
rect 17772 17380 17776 17436
rect 17776 17380 17832 17436
rect 17832 17380 17836 17436
rect 17772 17376 17836 17380
rect 17852 17436 17916 17440
rect 17852 17380 17856 17436
rect 17856 17380 17912 17436
rect 17912 17380 17916 17436
rect 17852 17376 17916 17380
rect 3372 17036 3436 17100
rect 2452 16960 2516 16964
rect 15148 17036 15212 17100
rect 2452 16904 2466 16960
rect 2466 16904 2516 16960
rect 2452 16900 2516 16904
rect 1952 16892 2016 16896
rect 1952 16836 1956 16892
rect 1956 16836 2012 16892
rect 2012 16836 2016 16892
rect 1952 16832 2016 16836
rect 2032 16892 2096 16896
rect 2032 16836 2036 16892
rect 2036 16836 2092 16892
rect 2092 16836 2096 16892
rect 2032 16832 2096 16836
rect 2112 16892 2176 16896
rect 2112 16836 2116 16892
rect 2116 16836 2172 16892
rect 2172 16836 2176 16892
rect 2112 16832 2176 16836
rect 2192 16892 2256 16896
rect 2192 16836 2196 16892
rect 2196 16836 2252 16892
rect 2252 16836 2256 16892
rect 2192 16832 2256 16836
rect 6952 16892 7016 16896
rect 6952 16836 6956 16892
rect 6956 16836 7012 16892
rect 7012 16836 7016 16892
rect 6952 16832 7016 16836
rect 7032 16892 7096 16896
rect 7032 16836 7036 16892
rect 7036 16836 7092 16892
rect 7092 16836 7096 16892
rect 7032 16832 7096 16836
rect 7112 16892 7176 16896
rect 7112 16836 7116 16892
rect 7116 16836 7172 16892
rect 7172 16836 7176 16892
rect 7112 16832 7176 16836
rect 7192 16892 7256 16896
rect 7192 16836 7196 16892
rect 7196 16836 7252 16892
rect 7252 16836 7256 16892
rect 7192 16832 7256 16836
rect 11952 16892 12016 16896
rect 11952 16836 11956 16892
rect 11956 16836 12012 16892
rect 12012 16836 12016 16892
rect 11952 16832 12016 16836
rect 12032 16892 12096 16896
rect 12032 16836 12036 16892
rect 12036 16836 12092 16892
rect 12092 16836 12096 16892
rect 12032 16832 12096 16836
rect 12112 16892 12176 16896
rect 12112 16836 12116 16892
rect 12116 16836 12172 16892
rect 12172 16836 12176 16892
rect 12112 16832 12176 16836
rect 12192 16892 12256 16896
rect 12192 16836 12196 16892
rect 12196 16836 12252 16892
rect 12252 16836 12256 16892
rect 12192 16832 12256 16836
rect 16952 16892 17016 16896
rect 16952 16836 16956 16892
rect 16956 16836 17012 16892
rect 17012 16836 17016 16892
rect 16952 16832 17016 16836
rect 17032 16892 17096 16896
rect 17032 16836 17036 16892
rect 17036 16836 17092 16892
rect 17092 16836 17096 16892
rect 17032 16832 17096 16836
rect 17112 16892 17176 16896
rect 17112 16836 17116 16892
rect 17116 16836 17172 16892
rect 17172 16836 17176 16892
rect 17112 16832 17176 16836
rect 17192 16892 17256 16896
rect 17192 16836 17196 16892
rect 17196 16836 17252 16892
rect 17252 16836 17256 16892
rect 17192 16832 17256 16836
rect 5396 16824 5460 16828
rect 5396 16768 5446 16824
rect 5446 16768 5460 16824
rect 5396 16764 5460 16768
rect 9076 16764 9140 16828
rect 13308 16764 13372 16828
rect 6316 16628 6380 16692
rect 16620 16492 16684 16556
rect 2612 16348 2676 16352
rect 2612 16292 2616 16348
rect 2616 16292 2672 16348
rect 2672 16292 2676 16348
rect 2612 16288 2676 16292
rect 2692 16348 2756 16352
rect 2692 16292 2696 16348
rect 2696 16292 2752 16348
rect 2752 16292 2756 16348
rect 2692 16288 2756 16292
rect 2772 16348 2836 16352
rect 2772 16292 2776 16348
rect 2776 16292 2832 16348
rect 2832 16292 2836 16348
rect 2772 16288 2836 16292
rect 2852 16348 2916 16352
rect 2852 16292 2856 16348
rect 2856 16292 2912 16348
rect 2912 16292 2916 16348
rect 2852 16288 2916 16292
rect 7612 16348 7676 16352
rect 7612 16292 7616 16348
rect 7616 16292 7672 16348
rect 7672 16292 7676 16348
rect 7612 16288 7676 16292
rect 7692 16348 7756 16352
rect 7692 16292 7696 16348
rect 7696 16292 7752 16348
rect 7752 16292 7756 16348
rect 7692 16288 7756 16292
rect 7772 16348 7836 16352
rect 7772 16292 7776 16348
rect 7776 16292 7832 16348
rect 7832 16292 7836 16348
rect 7772 16288 7836 16292
rect 7852 16348 7916 16352
rect 7852 16292 7856 16348
rect 7856 16292 7912 16348
rect 7912 16292 7916 16348
rect 7852 16288 7916 16292
rect 12612 16348 12676 16352
rect 12612 16292 12616 16348
rect 12616 16292 12672 16348
rect 12672 16292 12676 16348
rect 12612 16288 12676 16292
rect 12692 16348 12756 16352
rect 12692 16292 12696 16348
rect 12696 16292 12752 16348
rect 12752 16292 12756 16348
rect 12692 16288 12756 16292
rect 12772 16348 12836 16352
rect 12772 16292 12776 16348
rect 12776 16292 12832 16348
rect 12832 16292 12836 16348
rect 12772 16288 12836 16292
rect 12852 16348 12916 16352
rect 12852 16292 12856 16348
rect 12856 16292 12912 16348
rect 12912 16292 12916 16348
rect 12852 16288 12916 16292
rect 17612 16348 17676 16352
rect 17612 16292 17616 16348
rect 17616 16292 17672 16348
rect 17672 16292 17676 16348
rect 17612 16288 17676 16292
rect 17692 16348 17756 16352
rect 17692 16292 17696 16348
rect 17696 16292 17752 16348
rect 17752 16292 17756 16348
rect 17692 16288 17756 16292
rect 17772 16348 17836 16352
rect 17772 16292 17776 16348
rect 17776 16292 17832 16348
rect 17832 16292 17836 16348
rect 17772 16288 17836 16292
rect 17852 16348 17916 16352
rect 17852 16292 17856 16348
rect 17856 16292 17912 16348
rect 17912 16292 17916 16348
rect 17852 16288 17916 16292
rect 9444 16220 9508 16284
rect 10732 16220 10796 16284
rect 4292 15948 4356 16012
rect 10180 15812 10244 15876
rect 14228 15812 14292 15876
rect 1952 15804 2016 15808
rect 1952 15748 1956 15804
rect 1956 15748 2012 15804
rect 2012 15748 2016 15804
rect 1952 15744 2016 15748
rect 2032 15804 2096 15808
rect 2032 15748 2036 15804
rect 2036 15748 2092 15804
rect 2092 15748 2096 15804
rect 2032 15744 2096 15748
rect 2112 15804 2176 15808
rect 2112 15748 2116 15804
rect 2116 15748 2172 15804
rect 2172 15748 2176 15804
rect 2112 15744 2176 15748
rect 2192 15804 2256 15808
rect 2192 15748 2196 15804
rect 2196 15748 2252 15804
rect 2252 15748 2256 15804
rect 2192 15744 2256 15748
rect 6952 15804 7016 15808
rect 6952 15748 6956 15804
rect 6956 15748 7012 15804
rect 7012 15748 7016 15804
rect 6952 15744 7016 15748
rect 7032 15804 7096 15808
rect 7032 15748 7036 15804
rect 7036 15748 7092 15804
rect 7092 15748 7096 15804
rect 7032 15744 7096 15748
rect 7112 15804 7176 15808
rect 7112 15748 7116 15804
rect 7116 15748 7172 15804
rect 7172 15748 7176 15804
rect 7112 15744 7176 15748
rect 7192 15804 7256 15808
rect 7192 15748 7196 15804
rect 7196 15748 7252 15804
rect 7252 15748 7256 15804
rect 7192 15744 7256 15748
rect 11952 15804 12016 15808
rect 11952 15748 11956 15804
rect 11956 15748 12012 15804
rect 12012 15748 12016 15804
rect 11952 15744 12016 15748
rect 12032 15804 12096 15808
rect 12032 15748 12036 15804
rect 12036 15748 12092 15804
rect 12092 15748 12096 15804
rect 12032 15744 12096 15748
rect 12112 15804 12176 15808
rect 12112 15748 12116 15804
rect 12116 15748 12172 15804
rect 12172 15748 12176 15804
rect 12112 15744 12176 15748
rect 12192 15804 12256 15808
rect 12192 15748 12196 15804
rect 12196 15748 12252 15804
rect 12252 15748 12256 15804
rect 12192 15744 12256 15748
rect 16952 15804 17016 15808
rect 16952 15748 16956 15804
rect 16956 15748 17012 15804
rect 17012 15748 17016 15804
rect 16952 15744 17016 15748
rect 17032 15804 17096 15808
rect 17032 15748 17036 15804
rect 17036 15748 17092 15804
rect 17092 15748 17096 15804
rect 17032 15744 17096 15748
rect 17112 15804 17176 15808
rect 17112 15748 17116 15804
rect 17116 15748 17172 15804
rect 17172 15748 17176 15804
rect 17112 15744 17176 15748
rect 17192 15804 17256 15808
rect 17192 15748 17196 15804
rect 17196 15748 17252 15804
rect 17252 15748 17256 15804
rect 17192 15744 17256 15748
rect 9260 15404 9324 15468
rect 10916 15404 10980 15468
rect 18276 15404 18340 15468
rect 796 15268 860 15332
rect 4108 15268 4172 15332
rect 8708 15268 8772 15332
rect 2612 15260 2676 15264
rect 2612 15204 2616 15260
rect 2616 15204 2672 15260
rect 2672 15204 2676 15260
rect 2612 15200 2676 15204
rect 2692 15260 2756 15264
rect 2692 15204 2696 15260
rect 2696 15204 2752 15260
rect 2752 15204 2756 15260
rect 2692 15200 2756 15204
rect 2772 15260 2836 15264
rect 2772 15204 2776 15260
rect 2776 15204 2832 15260
rect 2832 15204 2836 15260
rect 2772 15200 2836 15204
rect 2852 15260 2916 15264
rect 2852 15204 2856 15260
rect 2856 15204 2912 15260
rect 2912 15204 2916 15260
rect 2852 15200 2916 15204
rect 7612 15260 7676 15264
rect 7612 15204 7616 15260
rect 7616 15204 7672 15260
rect 7672 15204 7676 15260
rect 7612 15200 7676 15204
rect 7692 15260 7756 15264
rect 7692 15204 7696 15260
rect 7696 15204 7752 15260
rect 7752 15204 7756 15260
rect 7692 15200 7756 15204
rect 7772 15260 7836 15264
rect 7772 15204 7776 15260
rect 7776 15204 7832 15260
rect 7832 15204 7836 15260
rect 7772 15200 7836 15204
rect 7852 15260 7916 15264
rect 7852 15204 7856 15260
rect 7856 15204 7912 15260
rect 7912 15204 7916 15260
rect 7852 15200 7916 15204
rect 12612 15260 12676 15264
rect 12612 15204 12616 15260
rect 12616 15204 12672 15260
rect 12672 15204 12676 15260
rect 12612 15200 12676 15204
rect 12692 15260 12756 15264
rect 12692 15204 12696 15260
rect 12696 15204 12752 15260
rect 12752 15204 12756 15260
rect 12692 15200 12756 15204
rect 12772 15260 12836 15264
rect 12772 15204 12776 15260
rect 12776 15204 12832 15260
rect 12832 15204 12836 15260
rect 12772 15200 12836 15204
rect 12852 15260 12916 15264
rect 12852 15204 12856 15260
rect 12856 15204 12912 15260
rect 12912 15204 12916 15260
rect 12852 15200 12916 15204
rect 17612 15260 17676 15264
rect 17612 15204 17616 15260
rect 17616 15204 17672 15260
rect 17672 15204 17676 15260
rect 17612 15200 17676 15204
rect 17692 15260 17756 15264
rect 17692 15204 17696 15260
rect 17696 15204 17752 15260
rect 17752 15204 17756 15260
rect 17692 15200 17756 15204
rect 17772 15260 17836 15264
rect 17772 15204 17776 15260
rect 17776 15204 17832 15260
rect 17832 15204 17836 15260
rect 17772 15200 17836 15204
rect 17852 15260 17916 15264
rect 17852 15204 17856 15260
rect 17856 15204 17912 15260
rect 17912 15204 17916 15260
rect 17852 15200 17916 15204
rect 7420 15132 7484 15196
rect 9628 15132 9692 15196
rect 8524 14996 8588 15060
rect 9812 15056 9876 15060
rect 9812 15000 9826 15056
rect 9826 15000 9876 15056
rect 9812 14996 9876 15000
rect 7420 14724 7484 14788
rect 13124 14724 13188 14788
rect 1952 14716 2016 14720
rect 1952 14660 1956 14716
rect 1956 14660 2012 14716
rect 2012 14660 2016 14716
rect 1952 14656 2016 14660
rect 2032 14716 2096 14720
rect 2032 14660 2036 14716
rect 2036 14660 2092 14716
rect 2092 14660 2096 14716
rect 2032 14656 2096 14660
rect 2112 14716 2176 14720
rect 2112 14660 2116 14716
rect 2116 14660 2172 14716
rect 2172 14660 2176 14716
rect 2112 14656 2176 14660
rect 2192 14716 2256 14720
rect 2192 14660 2196 14716
rect 2196 14660 2252 14716
rect 2252 14660 2256 14716
rect 2192 14656 2256 14660
rect 6952 14716 7016 14720
rect 6952 14660 6956 14716
rect 6956 14660 7012 14716
rect 7012 14660 7016 14716
rect 6952 14656 7016 14660
rect 7032 14716 7096 14720
rect 7032 14660 7036 14716
rect 7036 14660 7092 14716
rect 7092 14660 7096 14716
rect 7032 14656 7096 14660
rect 7112 14716 7176 14720
rect 7112 14660 7116 14716
rect 7116 14660 7172 14716
rect 7172 14660 7176 14716
rect 7112 14656 7176 14660
rect 7192 14716 7256 14720
rect 7192 14660 7196 14716
rect 7196 14660 7252 14716
rect 7252 14660 7256 14716
rect 7192 14656 7256 14660
rect 11952 14716 12016 14720
rect 11952 14660 11956 14716
rect 11956 14660 12012 14716
rect 12012 14660 12016 14716
rect 11952 14656 12016 14660
rect 12032 14716 12096 14720
rect 12032 14660 12036 14716
rect 12036 14660 12092 14716
rect 12092 14660 12096 14716
rect 12032 14656 12096 14660
rect 12112 14716 12176 14720
rect 12112 14660 12116 14716
rect 12116 14660 12172 14716
rect 12172 14660 12176 14716
rect 12112 14656 12176 14660
rect 12192 14716 12256 14720
rect 12192 14660 12196 14716
rect 12196 14660 12252 14716
rect 12252 14660 12256 14716
rect 12192 14656 12256 14660
rect 16952 14716 17016 14720
rect 16952 14660 16956 14716
rect 16956 14660 17012 14716
rect 17012 14660 17016 14716
rect 16952 14656 17016 14660
rect 17032 14716 17096 14720
rect 17032 14660 17036 14716
rect 17036 14660 17092 14716
rect 17092 14660 17096 14716
rect 17032 14656 17096 14660
rect 17112 14716 17176 14720
rect 17112 14660 17116 14716
rect 17116 14660 17172 14716
rect 17172 14660 17176 14716
rect 17112 14656 17176 14660
rect 17192 14716 17256 14720
rect 17192 14660 17196 14716
rect 17196 14660 17252 14716
rect 17252 14660 17256 14716
rect 17192 14656 17256 14660
rect 3740 14588 3804 14652
rect 7420 14588 7484 14652
rect 8340 14588 8404 14652
rect 15700 14588 15764 14652
rect 11652 14452 11716 14516
rect 2452 14180 2516 14244
rect 3924 14180 3988 14244
rect 2612 14172 2676 14176
rect 2612 14116 2616 14172
rect 2616 14116 2672 14172
rect 2672 14116 2676 14172
rect 2612 14112 2676 14116
rect 2692 14172 2756 14176
rect 2692 14116 2696 14172
rect 2696 14116 2752 14172
rect 2752 14116 2756 14172
rect 2692 14112 2756 14116
rect 2772 14172 2836 14176
rect 2772 14116 2776 14172
rect 2776 14116 2832 14172
rect 2832 14116 2836 14172
rect 2772 14112 2836 14116
rect 2852 14172 2916 14176
rect 2852 14116 2856 14172
rect 2856 14116 2912 14172
rect 2912 14116 2916 14172
rect 2852 14112 2916 14116
rect 5212 14044 5276 14108
rect 14964 14316 15028 14380
rect 7612 14172 7676 14176
rect 7612 14116 7616 14172
rect 7616 14116 7672 14172
rect 7672 14116 7676 14172
rect 7612 14112 7676 14116
rect 7692 14172 7756 14176
rect 7692 14116 7696 14172
rect 7696 14116 7752 14172
rect 7752 14116 7756 14172
rect 7692 14112 7756 14116
rect 7772 14172 7836 14176
rect 7772 14116 7776 14172
rect 7776 14116 7832 14172
rect 7832 14116 7836 14172
rect 7772 14112 7836 14116
rect 7852 14172 7916 14176
rect 7852 14116 7856 14172
rect 7856 14116 7912 14172
rect 7912 14116 7916 14172
rect 7852 14112 7916 14116
rect 12612 14172 12676 14176
rect 12612 14116 12616 14172
rect 12616 14116 12672 14172
rect 12672 14116 12676 14172
rect 12612 14112 12676 14116
rect 12692 14172 12756 14176
rect 12692 14116 12696 14172
rect 12696 14116 12752 14172
rect 12752 14116 12756 14172
rect 12692 14112 12756 14116
rect 12772 14172 12836 14176
rect 12772 14116 12776 14172
rect 12776 14116 12832 14172
rect 12832 14116 12836 14172
rect 12772 14112 12836 14116
rect 12852 14172 12916 14176
rect 12852 14116 12856 14172
rect 12856 14116 12912 14172
rect 12912 14116 12916 14172
rect 12852 14112 12916 14116
rect 17612 14172 17676 14176
rect 17612 14116 17616 14172
rect 17616 14116 17672 14172
rect 17672 14116 17676 14172
rect 17612 14112 17676 14116
rect 17692 14172 17756 14176
rect 17692 14116 17696 14172
rect 17696 14116 17752 14172
rect 17752 14116 17756 14172
rect 17692 14112 17756 14116
rect 17772 14172 17836 14176
rect 17772 14116 17776 14172
rect 17776 14116 17832 14172
rect 17832 14116 17836 14172
rect 17772 14112 17836 14116
rect 17852 14172 17916 14176
rect 17852 14116 17856 14172
rect 17856 14116 17912 14172
rect 17912 14116 17916 14172
rect 17852 14112 17916 14116
rect 18828 13908 18892 13972
rect 1164 13772 1228 13836
rect 6500 13832 6564 13836
rect 6500 13776 6514 13832
rect 6514 13776 6564 13832
rect 6500 13772 6564 13776
rect 3188 13636 3252 13700
rect 16620 13772 16684 13836
rect 8524 13636 8588 13700
rect 11468 13636 11532 13700
rect 1952 13628 2016 13632
rect 1952 13572 1956 13628
rect 1956 13572 2012 13628
rect 2012 13572 2016 13628
rect 1952 13568 2016 13572
rect 2032 13628 2096 13632
rect 2032 13572 2036 13628
rect 2036 13572 2092 13628
rect 2092 13572 2096 13628
rect 2032 13568 2096 13572
rect 2112 13628 2176 13632
rect 2112 13572 2116 13628
rect 2116 13572 2172 13628
rect 2172 13572 2176 13628
rect 2112 13568 2176 13572
rect 2192 13628 2256 13632
rect 2192 13572 2196 13628
rect 2196 13572 2252 13628
rect 2252 13572 2256 13628
rect 2192 13568 2256 13572
rect 6952 13628 7016 13632
rect 6952 13572 6956 13628
rect 6956 13572 7012 13628
rect 7012 13572 7016 13628
rect 6952 13568 7016 13572
rect 7032 13628 7096 13632
rect 7032 13572 7036 13628
rect 7036 13572 7092 13628
rect 7092 13572 7096 13628
rect 7032 13568 7096 13572
rect 7112 13628 7176 13632
rect 7112 13572 7116 13628
rect 7116 13572 7172 13628
rect 7172 13572 7176 13628
rect 7112 13568 7176 13572
rect 7192 13628 7256 13632
rect 7192 13572 7196 13628
rect 7196 13572 7252 13628
rect 7252 13572 7256 13628
rect 7192 13568 7256 13572
rect 11952 13628 12016 13632
rect 11952 13572 11956 13628
rect 11956 13572 12012 13628
rect 12012 13572 12016 13628
rect 11952 13568 12016 13572
rect 12032 13628 12096 13632
rect 12032 13572 12036 13628
rect 12036 13572 12092 13628
rect 12092 13572 12096 13628
rect 12032 13568 12096 13572
rect 12112 13628 12176 13632
rect 12112 13572 12116 13628
rect 12116 13572 12172 13628
rect 12172 13572 12176 13628
rect 12112 13568 12176 13572
rect 12192 13628 12256 13632
rect 12192 13572 12196 13628
rect 12196 13572 12252 13628
rect 12252 13572 12256 13628
rect 12192 13568 12256 13572
rect 16952 13628 17016 13632
rect 16952 13572 16956 13628
rect 16956 13572 17012 13628
rect 17012 13572 17016 13628
rect 16952 13568 17016 13572
rect 17032 13628 17096 13632
rect 17032 13572 17036 13628
rect 17036 13572 17092 13628
rect 17092 13572 17096 13628
rect 17032 13568 17096 13572
rect 17112 13628 17176 13632
rect 17112 13572 17116 13628
rect 17116 13572 17172 13628
rect 17172 13572 17176 13628
rect 17112 13568 17176 13572
rect 17192 13628 17256 13632
rect 17192 13572 17196 13628
rect 17196 13572 17252 13628
rect 17252 13572 17256 13628
rect 17192 13568 17256 13572
rect 1348 13364 1412 13428
rect 3004 13364 3068 13428
rect 5764 13500 5828 13564
rect 5948 13500 6012 13564
rect 6684 13500 6748 13564
rect 18644 13500 18708 13564
rect 4844 13364 4908 13428
rect 9996 13364 10060 13428
rect 10548 13364 10612 13428
rect 10364 13228 10428 13292
rect 11100 13228 11164 13292
rect 8524 13152 8588 13156
rect 8524 13096 8538 13152
rect 8538 13096 8588 13152
rect 8524 13092 8588 13096
rect 9076 13092 9140 13156
rect 2612 13084 2676 13088
rect 2612 13028 2616 13084
rect 2616 13028 2672 13084
rect 2672 13028 2676 13084
rect 2612 13024 2676 13028
rect 2692 13084 2756 13088
rect 2692 13028 2696 13084
rect 2696 13028 2752 13084
rect 2752 13028 2756 13084
rect 2692 13024 2756 13028
rect 2772 13084 2836 13088
rect 2772 13028 2776 13084
rect 2776 13028 2832 13084
rect 2832 13028 2836 13084
rect 2772 13024 2836 13028
rect 2852 13084 2916 13088
rect 2852 13028 2856 13084
rect 2856 13028 2912 13084
rect 2912 13028 2916 13084
rect 2852 13024 2916 13028
rect 7612 13084 7676 13088
rect 7612 13028 7616 13084
rect 7616 13028 7672 13084
rect 7672 13028 7676 13084
rect 7612 13024 7676 13028
rect 7692 13084 7756 13088
rect 7692 13028 7696 13084
rect 7696 13028 7752 13084
rect 7752 13028 7756 13084
rect 7692 13024 7756 13028
rect 7772 13084 7836 13088
rect 7772 13028 7776 13084
rect 7776 13028 7832 13084
rect 7832 13028 7836 13084
rect 7772 13024 7836 13028
rect 7852 13084 7916 13088
rect 7852 13028 7856 13084
rect 7856 13028 7912 13084
rect 7912 13028 7916 13084
rect 7852 13024 7916 13028
rect 4660 12956 4724 13020
rect 9076 12956 9140 13020
rect 9812 13092 9876 13156
rect 12612 13084 12676 13088
rect 12612 13028 12616 13084
rect 12616 13028 12672 13084
rect 12672 13028 12676 13084
rect 12612 13024 12676 13028
rect 12692 13084 12756 13088
rect 12692 13028 12696 13084
rect 12696 13028 12752 13084
rect 12752 13028 12756 13084
rect 12692 13024 12756 13028
rect 12772 13084 12836 13088
rect 12772 13028 12776 13084
rect 12776 13028 12832 13084
rect 12832 13028 12836 13084
rect 12772 13024 12836 13028
rect 12852 13084 12916 13088
rect 12852 13028 12856 13084
rect 12856 13028 12912 13084
rect 12912 13028 12916 13084
rect 12852 13024 12916 13028
rect 17612 13084 17676 13088
rect 17612 13028 17616 13084
rect 17616 13028 17672 13084
rect 17672 13028 17676 13084
rect 17612 13024 17676 13028
rect 17692 13084 17756 13088
rect 17692 13028 17696 13084
rect 17696 13028 17752 13084
rect 17752 13028 17756 13084
rect 17692 13024 17756 13028
rect 17772 13084 17836 13088
rect 17772 13028 17776 13084
rect 17776 13028 17832 13084
rect 17832 13028 17836 13084
rect 17772 13024 17836 13028
rect 17852 13084 17916 13088
rect 17852 13028 17856 13084
rect 17856 13028 17912 13084
rect 17912 13028 17916 13084
rect 17852 13024 17916 13028
rect 10548 12956 10612 13020
rect 19012 12820 19076 12884
rect 8892 12684 8956 12748
rect 9812 12744 9876 12748
rect 9812 12688 9826 12744
rect 9826 12688 9876 12744
rect 9812 12684 9876 12688
rect 10916 12548 10980 12612
rect 1952 12540 2016 12544
rect 1952 12484 1956 12540
rect 1956 12484 2012 12540
rect 2012 12484 2016 12540
rect 1952 12480 2016 12484
rect 2032 12540 2096 12544
rect 2032 12484 2036 12540
rect 2036 12484 2092 12540
rect 2092 12484 2096 12540
rect 2032 12480 2096 12484
rect 2112 12540 2176 12544
rect 2112 12484 2116 12540
rect 2116 12484 2172 12540
rect 2172 12484 2176 12540
rect 2112 12480 2176 12484
rect 2192 12540 2256 12544
rect 2192 12484 2196 12540
rect 2196 12484 2252 12540
rect 2252 12484 2256 12540
rect 2192 12480 2256 12484
rect 6952 12540 7016 12544
rect 6952 12484 6956 12540
rect 6956 12484 7012 12540
rect 7012 12484 7016 12540
rect 6952 12480 7016 12484
rect 7032 12540 7096 12544
rect 7032 12484 7036 12540
rect 7036 12484 7092 12540
rect 7092 12484 7096 12540
rect 7032 12480 7096 12484
rect 7112 12540 7176 12544
rect 7112 12484 7116 12540
rect 7116 12484 7172 12540
rect 7172 12484 7176 12540
rect 7112 12480 7176 12484
rect 7192 12540 7256 12544
rect 7192 12484 7196 12540
rect 7196 12484 7252 12540
rect 7252 12484 7256 12540
rect 7192 12480 7256 12484
rect 11952 12540 12016 12544
rect 11952 12484 11956 12540
rect 11956 12484 12012 12540
rect 12012 12484 12016 12540
rect 11952 12480 12016 12484
rect 12032 12540 12096 12544
rect 12032 12484 12036 12540
rect 12036 12484 12092 12540
rect 12092 12484 12096 12540
rect 12032 12480 12096 12484
rect 12112 12540 12176 12544
rect 12112 12484 12116 12540
rect 12116 12484 12172 12540
rect 12172 12484 12176 12540
rect 12112 12480 12176 12484
rect 12192 12540 12256 12544
rect 12192 12484 12196 12540
rect 12196 12484 12252 12540
rect 12252 12484 12256 12540
rect 12192 12480 12256 12484
rect 16952 12540 17016 12544
rect 16952 12484 16956 12540
rect 16956 12484 17012 12540
rect 17012 12484 17016 12540
rect 16952 12480 17016 12484
rect 17032 12540 17096 12544
rect 17032 12484 17036 12540
rect 17036 12484 17092 12540
rect 17092 12484 17096 12540
rect 17032 12480 17096 12484
rect 17112 12540 17176 12544
rect 17112 12484 17116 12540
rect 17116 12484 17172 12540
rect 17172 12484 17176 12540
rect 17112 12480 17176 12484
rect 17192 12540 17256 12544
rect 17192 12484 17196 12540
rect 17196 12484 17252 12540
rect 17252 12484 17256 12540
rect 17192 12480 17256 12484
rect 5028 12276 5092 12340
rect 5764 12336 5828 12340
rect 5764 12280 5814 12336
rect 5814 12280 5828 12336
rect 5764 12276 5828 12280
rect 8156 12004 8220 12068
rect 9260 12004 9324 12068
rect 11284 12140 11348 12204
rect 12388 12140 12452 12204
rect 13308 12140 13372 12204
rect 2612 11996 2676 12000
rect 2612 11940 2616 11996
rect 2616 11940 2672 11996
rect 2672 11940 2676 11996
rect 2612 11936 2676 11940
rect 2692 11996 2756 12000
rect 2692 11940 2696 11996
rect 2696 11940 2752 11996
rect 2752 11940 2756 11996
rect 2692 11936 2756 11940
rect 2772 11996 2836 12000
rect 2772 11940 2776 11996
rect 2776 11940 2832 11996
rect 2832 11940 2836 11996
rect 2772 11936 2836 11940
rect 2852 11996 2916 12000
rect 2852 11940 2856 11996
rect 2856 11940 2912 11996
rect 2912 11940 2916 11996
rect 2852 11936 2916 11940
rect 7612 11996 7676 12000
rect 7612 11940 7616 11996
rect 7616 11940 7672 11996
rect 7672 11940 7676 11996
rect 7612 11936 7676 11940
rect 7692 11996 7756 12000
rect 7692 11940 7696 11996
rect 7696 11940 7752 11996
rect 7752 11940 7756 11996
rect 7692 11936 7756 11940
rect 7772 11996 7836 12000
rect 7772 11940 7776 11996
rect 7776 11940 7832 11996
rect 7832 11940 7836 11996
rect 7772 11936 7836 11940
rect 7852 11996 7916 12000
rect 7852 11940 7856 11996
rect 7856 11940 7912 11996
rect 7912 11940 7916 11996
rect 7852 11936 7916 11940
rect 12612 11996 12676 12000
rect 12612 11940 12616 11996
rect 12616 11940 12672 11996
rect 12672 11940 12676 11996
rect 12612 11936 12676 11940
rect 12692 11996 12756 12000
rect 12692 11940 12696 11996
rect 12696 11940 12752 11996
rect 12752 11940 12756 11996
rect 12692 11936 12756 11940
rect 12772 11996 12836 12000
rect 12772 11940 12776 11996
rect 12776 11940 12832 11996
rect 12832 11940 12836 11996
rect 12772 11936 12836 11940
rect 12852 11996 12916 12000
rect 12852 11940 12856 11996
rect 12856 11940 12912 11996
rect 12912 11940 12916 11996
rect 12852 11936 12916 11940
rect 5028 11732 5092 11796
rect 15148 12276 15212 12340
rect 13676 12140 13740 12204
rect 15148 12140 15212 12204
rect 18460 12140 18524 12204
rect 17612 11996 17676 12000
rect 17612 11940 17616 11996
rect 17616 11940 17672 11996
rect 17672 11940 17676 11996
rect 17612 11936 17676 11940
rect 17692 11996 17756 12000
rect 17692 11940 17696 11996
rect 17696 11940 17752 11996
rect 17752 11940 17756 11996
rect 17692 11936 17756 11940
rect 17772 11996 17836 12000
rect 17772 11940 17776 11996
rect 17776 11940 17832 11996
rect 17832 11940 17836 11996
rect 17772 11936 17836 11940
rect 17852 11996 17916 12000
rect 17852 11940 17856 11996
rect 17856 11940 17912 11996
rect 17912 11940 17916 11996
rect 17852 11936 17916 11940
rect 16252 11868 16316 11932
rect 10180 11732 10244 11796
rect 10916 11792 10980 11796
rect 10916 11736 10930 11792
rect 10930 11736 10980 11792
rect 10916 11732 10980 11736
rect 2452 11460 2516 11524
rect 1952 11452 2016 11456
rect 1952 11396 1956 11452
rect 1956 11396 2012 11452
rect 2012 11396 2016 11452
rect 1952 11392 2016 11396
rect 2032 11452 2096 11456
rect 2032 11396 2036 11452
rect 2036 11396 2092 11452
rect 2092 11396 2096 11452
rect 2032 11392 2096 11396
rect 2112 11452 2176 11456
rect 2112 11396 2116 11452
rect 2116 11396 2172 11452
rect 2172 11396 2176 11452
rect 2112 11392 2176 11396
rect 2192 11452 2256 11456
rect 2192 11396 2196 11452
rect 2196 11396 2252 11452
rect 2252 11396 2256 11452
rect 2192 11392 2256 11396
rect 6952 11452 7016 11456
rect 6952 11396 6956 11452
rect 6956 11396 7012 11452
rect 7012 11396 7016 11452
rect 6952 11392 7016 11396
rect 7032 11452 7096 11456
rect 7032 11396 7036 11452
rect 7036 11396 7092 11452
rect 7092 11396 7096 11452
rect 7032 11392 7096 11396
rect 7112 11452 7176 11456
rect 7112 11396 7116 11452
rect 7116 11396 7172 11452
rect 7172 11396 7176 11452
rect 7112 11392 7176 11396
rect 7192 11452 7256 11456
rect 7192 11396 7196 11452
rect 7196 11396 7252 11452
rect 7252 11396 7256 11452
rect 7192 11392 7256 11396
rect 4476 11384 4540 11388
rect 4476 11328 4490 11384
rect 4490 11328 4540 11384
rect 4476 11324 4540 11328
rect 8340 11324 8404 11388
rect 9260 11384 9324 11388
rect 9260 11328 9274 11384
rect 9274 11328 9324 11384
rect 9260 11324 9324 11328
rect 9628 11324 9692 11388
rect 4660 11248 4724 11252
rect 4660 11192 4674 11248
rect 4674 11192 4724 11248
rect 4660 11188 4724 11192
rect 5580 11188 5644 11252
rect 10732 11188 10796 11252
rect 14044 11460 14108 11524
rect 14780 11520 14844 11524
rect 14780 11464 14830 11520
rect 14830 11464 14844 11520
rect 14780 11460 14844 11464
rect 11952 11452 12016 11456
rect 11952 11396 11956 11452
rect 11956 11396 12012 11452
rect 12012 11396 12016 11452
rect 11952 11392 12016 11396
rect 12032 11452 12096 11456
rect 12032 11396 12036 11452
rect 12036 11396 12092 11452
rect 12092 11396 12096 11452
rect 12032 11392 12096 11396
rect 12112 11452 12176 11456
rect 12112 11396 12116 11452
rect 12116 11396 12172 11452
rect 12172 11396 12176 11452
rect 12112 11392 12176 11396
rect 12192 11452 12256 11456
rect 12192 11396 12196 11452
rect 12196 11396 12252 11452
rect 12252 11396 12256 11452
rect 12192 11392 12256 11396
rect 16952 11452 17016 11456
rect 16952 11396 16956 11452
rect 16956 11396 17012 11452
rect 17012 11396 17016 11452
rect 16952 11392 17016 11396
rect 17032 11452 17096 11456
rect 17032 11396 17036 11452
rect 17036 11396 17092 11452
rect 17092 11396 17096 11452
rect 17032 11392 17096 11396
rect 17112 11452 17176 11456
rect 17112 11396 17116 11452
rect 17116 11396 17172 11452
rect 17172 11396 17176 11452
rect 17112 11392 17176 11396
rect 17192 11452 17256 11456
rect 17192 11396 17196 11452
rect 17196 11396 17252 11452
rect 17252 11396 17256 11452
rect 17192 11392 17256 11396
rect 16252 11324 16316 11388
rect 13860 11112 13924 11116
rect 13860 11056 13874 11112
rect 13874 11056 13924 11112
rect 3188 10916 3252 10980
rect 2612 10908 2676 10912
rect 2612 10852 2616 10908
rect 2616 10852 2672 10908
rect 2672 10852 2676 10908
rect 2612 10848 2676 10852
rect 2692 10908 2756 10912
rect 2692 10852 2696 10908
rect 2696 10852 2752 10908
rect 2752 10852 2756 10908
rect 2692 10848 2756 10852
rect 2772 10908 2836 10912
rect 2772 10852 2776 10908
rect 2776 10852 2832 10908
rect 2832 10852 2836 10908
rect 2772 10848 2836 10852
rect 2852 10908 2916 10912
rect 2852 10852 2856 10908
rect 2856 10852 2912 10908
rect 2912 10852 2916 10908
rect 2852 10848 2916 10852
rect 3556 10780 3620 10844
rect 4108 10780 4172 10844
rect 4292 10780 4356 10844
rect 5396 10780 5460 10844
rect 6316 10644 6380 10708
rect 7420 10916 7484 10980
rect 13860 11052 13924 11056
rect 15884 11052 15948 11116
rect 14596 10916 14660 10980
rect 15516 10916 15580 10980
rect 7612 10908 7676 10912
rect 7612 10852 7616 10908
rect 7616 10852 7672 10908
rect 7672 10852 7676 10908
rect 7612 10848 7676 10852
rect 7692 10908 7756 10912
rect 7692 10852 7696 10908
rect 7696 10852 7752 10908
rect 7752 10852 7756 10908
rect 7692 10848 7756 10852
rect 7772 10908 7836 10912
rect 7772 10852 7776 10908
rect 7776 10852 7832 10908
rect 7832 10852 7836 10908
rect 7772 10848 7836 10852
rect 7852 10908 7916 10912
rect 7852 10852 7856 10908
rect 7856 10852 7912 10908
rect 7912 10852 7916 10908
rect 7852 10848 7916 10852
rect 12612 10908 12676 10912
rect 12612 10852 12616 10908
rect 12616 10852 12672 10908
rect 12672 10852 12676 10908
rect 12612 10848 12676 10852
rect 12692 10908 12756 10912
rect 12692 10852 12696 10908
rect 12696 10852 12752 10908
rect 12752 10852 12756 10908
rect 12692 10848 12756 10852
rect 12772 10908 12836 10912
rect 12772 10852 12776 10908
rect 12776 10852 12832 10908
rect 12832 10852 12836 10908
rect 12772 10848 12836 10852
rect 12852 10908 12916 10912
rect 12852 10852 12856 10908
rect 12856 10852 12912 10908
rect 12912 10852 12916 10908
rect 12852 10848 12916 10852
rect 17612 10908 17676 10912
rect 17612 10852 17616 10908
rect 17616 10852 17672 10908
rect 17672 10852 17676 10908
rect 17612 10848 17676 10852
rect 17692 10908 17756 10912
rect 17692 10852 17696 10908
rect 17696 10852 17752 10908
rect 17752 10852 17756 10908
rect 17692 10848 17756 10852
rect 17772 10908 17836 10912
rect 17772 10852 17776 10908
rect 17776 10852 17832 10908
rect 17832 10852 17836 10908
rect 17772 10848 17836 10852
rect 17852 10908 17916 10912
rect 17852 10852 17856 10908
rect 17856 10852 17912 10908
rect 17912 10852 17916 10908
rect 17852 10848 17916 10852
rect 7420 10780 7484 10844
rect 10732 10780 10796 10844
rect 11284 10780 11348 10844
rect 15332 10840 15396 10844
rect 15332 10784 15346 10840
rect 15346 10784 15396 10840
rect 15332 10780 15396 10784
rect 15884 10840 15948 10844
rect 15884 10784 15934 10840
rect 15934 10784 15948 10840
rect 15884 10780 15948 10784
rect 3556 10372 3620 10436
rect 3740 10372 3804 10436
rect 6316 10508 6380 10572
rect 9444 10508 9508 10572
rect 11100 10644 11164 10708
rect 1952 10364 2016 10368
rect 1952 10308 1956 10364
rect 1956 10308 2012 10364
rect 2012 10308 2016 10364
rect 1952 10304 2016 10308
rect 2032 10364 2096 10368
rect 2032 10308 2036 10364
rect 2036 10308 2092 10364
rect 2092 10308 2096 10364
rect 2032 10304 2096 10308
rect 2112 10364 2176 10368
rect 2112 10308 2116 10364
rect 2116 10308 2172 10364
rect 2172 10308 2176 10364
rect 2112 10304 2176 10308
rect 2192 10364 2256 10368
rect 2192 10308 2196 10364
rect 2196 10308 2252 10364
rect 2252 10308 2256 10364
rect 2192 10304 2256 10308
rect 6952 10364 7016 10368
rect 6952 10308 6956 10364
rect 6956 10308 7012 10364
rect 7012 10308 7016 10364
rect 6952 10304 7016 10308
rect 7032 10364 7096 10368
rect 7032 10308 7036 10364
rect 7036 10308 7092 10364
rect 7092 10308 7096 10364
rect 7032 10304 7096 10308
rect 7112 10364 7176 10368
rect 7112 10308 7116 10364
rect 7116 10308 7172 10364
rect 7172 10308 7176 10364
rect 7112 10304 7176 10308
rect 7192 10364 7256 10368
rect 7192 10308 7196 10364
rect 7196 10308 7252 10364
rect 7252 10308 7256 10364
rect 7192 10304 7256 10308
rect 11952 10364 12016 10368
rect 11952 10308 11956 10364
rect 11956 10308 12012 10364
rect 12012 10308 12016 10364
rect 11952 10304 12016 10308
rect 12032 10364 12096 10368
rect 12032 10308 12036 10364
rect 12036 10308 12092 10364
rect 12092 10308 12096 10364
rect 12032 10304 12096 10308
rect 12112 10364 12176 10368
rect 12112 10308 12116 10364
rect 12116 10308 12172 10364
rect 12172 10308 12176 10364
rect 12112 10304 12176 10308
rect 12192 10364 12256 10368
rect 12192 10308 12196 10364
rect 12196 10308 12252 10364
rect 12252 10308 12256 10364
rect 12192 10304 12256 10308
rect 16952 10364 17016 10368
rect 16952 10308 16956 10364
rect 16956 10308 17012 10364
rect 17012 10308 17016 10364
rect 16952 10304 17016 10308
rect 17032 10364 17096 10368
rect 17032 10308 17036 10364
rect 17036 10308 17092 10364
rect 17092 10308 17096 10364
rect 17032 10304 17096 10308
rect 17112 10364 17176 10368
rect 17112 10308 17116 10364
rect 17116 10308 17172 10364
rect 17172 10308 17176 10364
rect 17112 10304 17176 10308
rect 17192 10364 17256 10368
rect 17192 10308 17196 10364
rect 17196 10308 17252 10364
rect 17252 10308 17256 10364
rect 17192 10304 17256 10308
rect 3188 10100 3252 10164
rect 5764 10236 5828 10300
rect 9444 10296 9508 10300
rect 9444 10240 9494 10296
rect 9494 10240 9508 10296
rect 9444 10236 9508 10240
rect 9628 10236 9692 10300
rect 10364 10236 10428 10300
rect 13492 10236 13556 10300
rect 15516 10100 15580 10164
rect 19380 10100 19444 10164
rect 3004 9828 3068 9892
rect 4292 10024 4356 10028
rect 4292 9968 4342 10024
rect 4342 9968 4356 10024
rect 4292 9964 4356 9968
rect 5580 9964 5644 10028
rect 2612 9820 2676 9824
rect 2612 9764 2616 9820
rect 2616 9764 2672 9820
rect 2672 9764 2676 9820
rect 2612 9760 2676 9764
rect 2692 9820 2756 9824
rect 2692 9764 2696 9820
rect 2696 9764 2752 9820
rect 2752 9764 2756 9820
rect 2692 9760 2756 9764
rect 2772 9820 2836 9824
rect 2772 9764 2776 9820
rect 2776 9764 2832 9820
rect 2832 9764 2836 9820
rect 2772 9760 2836 9764
rect 2852 9820 2916 9824
rect 2852 9764 2856 9820
rect 2856 9764 2912 9820
rect 2912 9764 2916 9820
rect 2852 9760 2916 9764
rect 3372 9556 3436 9620
rect 5028 9556 5092 9620
rect 6316 9692 6380 9756
rect 6316 9556 6380 9620
rect 13308 9828 13372 9892
rect 13860 9828 13924 9892
rect 15884 9828 15948 9892
rect 16436 9828 16500 9892
rect 7612 9820 7676 9824
rect 7612 9764 7616 9820
rect 7616 9764 7672 9820
rect 7672 9764 7676 9820
rect 7612 9760 7676 9764
rect 7692 9820 7756 9824
rect 7692 9764 7696 9820
rect 7696 9764 7752 9820
rect 7752 9764 7756 9820
rect 7692 9760 7756 9764
rect 7772 9820 7836 9824
rect 7772 9764 7776 9820
rect 7776 9764 7832 9820
rect 7832 9764 7836 9820
rect 7772 9760 7836 9764
rect 7852 9820 7916 9824
rect 7852 9764 7856 9820
rect 7856 9764 7912 9820
rect 7912 9764 7916 9820
rect 7852 9760 7916 9764
rect 12612 9820 12676 9824
rect 12612 9764 12616 9820
rect 12616 9764 12672 9820
rect 12672 9764 12676 9820
rect 12612 9760 12676 9764
rect 12692 9820 12756 9824
rect 12692 9764 12696 9820
rect 12696 9764 12752 9820
rect 12752 9764 12756 9820
rect 12692 9760 12756 9764
rect 12772 9820 12836 9824
rect 12772 9764 12776 9820
rect 12776 9764 12832 9820
rect 12832 9764 12836 9820
rect 12772 9760 12836 9764
rect 12852 9820 12916 9824
rect 12852 9764 12856 9820
rect 12856 9764 12912 9820
rect 12912 9764 12916 9820
rect 12852 9760 12916 9764
rect 17612 9820 17676 9824
rect 17612 9764 17616 9820
rect 17616 9764 17672 9820
rect 17672 9764 17676 9820
rect 17612 9760 17676 9764
rect 17692 9820 17756 9824
rect 17692 9764 17696 9820
rect 17696 9764 17752 9820
rect 17752 9764 17756 9820
rect 17692 9760 17756 9764
rect 17772 9820 17836 9824
rect 17772 9764 17776 9820
rect 17776 9764 17832 9820
rect 17832 9764 17836 9820
rect 17772 9760 17836 9764
rect 17852 9820 17916 9824
rect 17852 9764 17856 9820
rect 17856 9764 17912 9820
rect 17912 9764 17916 9820
rect 17852 9760 17916 9764
rect 9996 9692 10060 9756
rect 12388 9692 12452 9756
rect 13492 9692 13556 9756
rect 16068 9692 16132 9756
rect 18092 9692 18156 9756
rect 1716 9420 1780 9484
rect 2452 9420 2516 9484
rect 3188 9420 3252 9484
rect 5580 9420 5644 9484
rect 5764 9420 5828 9484
rect 16252 9556 16316 9620
rect 16804 9556 16868 9620
rect 3188 9284 3252 9348
rect 5028 9284 5092 9348
rect 5212 9284 5276 9348
rect 9076 9420 9140 9484
rect 14228 9344 14292 9348
rect 14228 9288 14278 9344
rect 14278 9288 14292 9344
rect 1952 9276 2016 9280
rect 1952 9220 1956 9276
rect 1956 9220 2012 9276
rect 2012 9220 2016 9276
rect 1952 9216 2016 9220
rect 2032 9276 2096 9280
rect 2032 9220 2036 9276
rect 2036 9220 2092 9276
rect 2092 9220 2096 9276
rect 2032 9216 2096 9220
rect 2112 9276 2176 9280
rect 2112 9220 2116 9276
rect 2116 9220 2172 9276
rect 2172 9220 2176 9276
rect 2112 9216 2176 9220
rect 2192 9276 2256 9280
rect 2192 9220 2196 9276
rect 2196 9220 2252 9276
rect 2252 9220 2256 9276
rect 2192 9216 2256 9220
rect 6952 9276 7016 9280
rect 6952 9220 6956 9276
rect 6956 9220 7012 9276
rect 7012 9220 7016 9276
rect 6952 9216 7016 9220
rect 7032 9276 7096 9280
rect 7032 9220 7036 9276
rect 7036 9220 7092 9276
rect 7092 9220 7096 9276
rect 7032 9216 7096 9220
rect 7112 9276 7176 9280
rect 7112 9220 7116 9276
rect 7116 9220 7172 9276
rect 7172 9220 7176 9276
rect 7112 9216 7176 9220
rect 7192 9276 7256 9280
rect 7192 9220 7196 9276
rect 7196 9220 7252 9276
rect 7252 9220 7256 9276
rect 7192 9216 7256 9220
rect 796 9072 860 9076
rect 796 9016 810 9072
rect 810 9016 860 9072
rect 796 9012 860 9016
rect 4660 9148 4724 9212
rect 6316 9148 6380 9212
rect 8156 9148 8220 9212
rect 10180 9148 10244 9212
rect 4108 9012 4172 9076
rect 8892 9012 8956 9076
rect 10732 9012 10796 9076
rect 11284 9012 11348 9076
rect 14228 9284 14292 9288
rect 14412 9344 14476 9348
rect 14412 9288 14462 9344
rect 14462 9288 14476 9344
rect 14412 9284 14476 9288
rect 11952 9276 12016 9280
rect 11952 9220 11956 9276
rect 11956 9220 12012 9276
rect 12012 9220 12016 9276
rect 11952 9216 12016 9220
rect 12032 9276 12096 9280
rect 12032 9220 12036 9276
rect 12036 9220 12092 9276
rect 12092 9220 12096 9276
rect 12032 9216 12096 9220
rect 12112 9276 12176 9280
rect 12112 9220 12116 9276
rect 12116 9220 12172 9276
rect 12172 9220 12176 9276
rect 12112 9216 12176 9220
rect 12192 9276 12256 9280
rect 12192 9220 12196 9276
rect 12196 9220 12252 9276
rect 12252 9220 12256 9276
rect 12192 9216 12256 9220
rect 16252 9420 16316 9484
rect 16952 9276 17016 9280
rect 16952 9220 16956 9276
rect 16956 9220 17012 9276
rect 17012 9220 17016 9276
rect 16952 9216 17016 9220
rect 17032 9276 17096 9280
rect 17032 9220 17036 9276
rect 17036 9220 17092 9276
rect 17092 9220 17096 9276
rect 17032 9216 17096 9220
rect 17112 9276 17176 9280
rect 17112 9220 17116 9276
rect 17116 9220 17172 9276
rect 17172 9220 17176 9276
rect 17112 9216 17176 9220
rect 17192 9276 17256 9280
rect 17192 9220 17196 9276
rect 17196 9220 17252 9276
rect 17252 9220 17256 9276
rect 17192 9216 17256 9220
rect 4660 8876 4724 8940
rect 6316 8876 6380 8940
rect 2612 8732 2676 8736
rect 2612 8676 2616 8732
rect 2616 8676 2672 8732
rect 2672 8676 2676 8732
rect 2612 8672 2676 8676
rect 2692 8732 2756 8736
rect 2692 8676 2696 8732
rect 2696 8676 2752 8732
rect 2752 8676 2756 8732
rect 2692 8672 2756 8676
rect 2772 8732 2836 8736
rect 2772 8676 2776 8732
rect 2776 8676 2832 8732
rect 2832 8676 2836 8732
rect 2772 8672 2836 8676
rect 2852 8732 2916 8736
rect 2852 8676 2856 8732
rect 2856 8676 2912 8732
rect 2912 8676 2916 8732
rect 2852 8672 2916 8676
rect 1532 8604 1596 8668
rect 1348 8468 1412 8532
rect 3004 8468 3068 8532
rect 3372 8332 3436 8396
rect 5396 8604 5460 8668
rect 6684 8740 6748 8804
rect 8892 8740 8956 8804
rect 7612 8732 7676 8736
rect 7612 8676 7616 8732
rect 7616 8676 7672 8732
rect 7672 8676 7676 8732
rect 7612 8672 7676 8676
rect 7692 8732 7756 8736
rect 7692 8676 7696 8732
rect 7696 8676 7752 8732
rect 7752 8676 7756 8732
rect 7692 8672 7756 8676
rect 7772 8732 7836 8736
rect 7772 8676 7776 8732
rect 7776 8676 7832 8732
rect 7832 8676 7836 8732
rect 7772 8672 7836 8676
rect 7852 8732 7916 8736
rect 7852 8676 7856 8732
rect 7856 8676 7912 8732
rect 7912 8676 7916 8732
rect 7852 8672 7916 8676
rect 12612 8732 12676 8736
rect 12612 8676 12616 8732
rect 12616 8676 12672 8732
rect 12672 8676 12676 8732
rect 12612 8672 12676 8676
rect 12692 8732 12756 8736
rect 12692 8676 12696 8732
rect 12696 8676 12752 8732
rect 12752 8676 12756 8732
rect 12692 8672 12756 8676
rect 12772 8732 12836 8736
rect 12772 8676 12776 8732
rect 12776 8676 12832 8732
rect 12832 8676 12836 8732
rect 12772 8672 12836 8676
rect 12852 8732 12916 8736
rect 12852 8676 12856 8732
rect 12856 8676 12912 8732
rect 12912 8676 12916 8732
rect 12852 8672 12916 8676
rect 17612 8732 17676 8736
rect 17612 8676 17616 8732
rect 17616 8676 17672 8732
rect 17672 8676 17676 8732
rect 17612 8672 17676 8676
rect 17692 8732 17756 8736
rect 17692 8676 17696 8732
rect 17696 8676 17752 8732
rect 17752 8676 17756 8732
rect 17692 8672 17756 8676
rect 17772 8732 17836 8736
rect 17772 8676 17776 8732
rect 17776 8676 17832 8732
rect 17832 8676 17836 8732
rect 17772 8672 17836 8676
rect 17852 8732 17916 8736
rect 17852 8676 17856 8732
rect 17856 8676 17912 8732
rect 17912 8676 17916 8732
rect 17852 8672 17916 8676
rect 9996 8468 10060 8532
rect 5396 8332 5460 8396
rect 13308 8332 13372 8396
rect 4108 8196 4172 8260
rect 1952 8188 2016 8192
rect 1952 8132 1956 8188
rect 1956 8132 2012 8188
rect 2012 8132 2016 8188
rect 1952 8128 2016 8132
rect 2032 8188 2096 8192
rect 2032 8132 2036 8188
rect 2036 8132 2092 8188
rect 2092 8132 2096 8188
rect 2032 8128 2096 8132
rect 2112 8188 2176 8192
rect 2112 8132 2116 8188
rect 2116 8132 2172 8188
rect 2172 8132 2176 8188
rect 2112 8128 2176 8132
rect 2192 8188 2256 8192
rect 2192 8132 2196 8188
rect 2196 8132 2252 8188
rect 2252 8132 2256 8188
rect 2192 8128 2256 8132
rect 3740 8060 3804 8124
rect 5948 8060 6012 8124
rect 6684 8256 6748 8260
rect 6684 8200 6698 8256
rect 6698 8200 6748 8256
rect 6684 8196 6748 8200
rect 7420 8196 7484 8260
rect 8340 8196 8404 8260
rect 10732 8196 10796 8260
rect 6952 8188 7016 8192
rect 6952 8132 6956 8188
rect 6956 8132 7012 8188
rect 7012 8132 7016 8188
rect 6952 8128 7016 8132
rect 7032 8188 7096 8192
rect 7032 8132 7036 8188
rect 7036 8132 7092 8188
rect 7092 8132 7096 8188
rect 7032 8128 7096 8132
rect 7112 8188 7176 8192
rect 7112 8132 7116 8188
rect 7116 8132 7172 8188
rect 7172 8132 7176 8188
rect 7112 8128 7176 8132
rect 7192 8188 7256 8192
rect 7192 8132 7196 8188
rect 7196 8132 7252 8188
rect 7252 8132 7256 8188
rect 7192 8128 7256 8132
rect 11952 8188 12016 8192
rect 11952 8132 11956 8188
rect 11956 8132 12012 8188
rect 12012 8132 12016 8188
rect 11952 8128 12016 8132
rect 12032 8188 12096 8192
rect 12032 8132 12036 8188
rect 12036 8132 12092 8188
rect 12092 8132 12096 8188
rect 12032 8128 12096 8132
rect 12112 8188 12176 8192
rect 12112 8132 12116 8188
rect 12116 8132 12172 8188
rect 12172 8132 12176 8188
rect 12112 8128 12176 8132
rect 12192 8188 12256 8192
rect 12192 8132 12196 8188
rect 12196 8132 12252 8188
rect 12252 8132 12256 8188
rect 12192 8128 12256 8132
rect 9444 8060 9508 8124
rect 16952 8188 17016 8192
rect 16952 8132 16956 8188
rect 16956 8132 17012 8188
rect 17012 8132 17016 8188
rect 16952 8128 17016 8132
rect 17032 8188 17096 8192
rect 17032 8132 17036 8188
rect 17036 8132 17092 8188
rect 17092 8132 17096 8188
rect 17032 8128 17096 8132
rect 17112 8188 17176 8192
rect 17112 8132 17116 8188
rect 17116 8132 17172 8188
rect 17172 8132 17176 8188
rect 17112 8128 17176 8132
rect 17192 8188 17256 8192
rect 17192 8132 17196 8188
rect 17196 8132 17252 8188
rect 17252 8132 17256 8188
rect 17192 8128 17256 8132
rect 14596 8060 14660 8124
rect 3556 7924 3620 7988
rect 4660 7788 4724 7852
rect 8156 7984 8220 7988
rect 8156 7928 8170 7984
rect 8170 7928 8220 7984
rect 8156 7924 8220 7928
rect 5028 7652 5092 7716
rect 8340 7788 8404 7852
rect 15700 7924 15764 7988
rect 11100 7652 11164 7716
rect 11468 7652 11532 7716
rect 2612 7644 2676 7648
rect 2612 7588 2616 7644
rect 2616 7588 2672 7644
rect 2672 7588 2676 7644
rect 2612 7584 2676 7588
rect 2692 7644 2756 7648
rect 2692 7588 2696 7644
rect 2696 7588 2752 7644
rect 2752 7588 2756 7644
rect 2692 7584 2756 7588
rect 2772 7644 2836 7648
rect 2772 7588 2776 7644
rect 2776 7588 2832 7644
rect 2832 7588 2836 7644
rect 2772 7584 2836 7588
rect 2852 7644 2916 7648
rect 2852 7588 2856 7644
rect 2856 7588 2912 7644
rect 2912 7588 2916 7644
rect 2852 7584 2916 7588
rect 7612 7644 7676 7648
rect 7612 7588 7616 7644
rect 7616 7588 7672 7644
rect 7672 7588 7676 7644
rect 7612 7584 7676 7588
rect 7692 7644 7756 7648
rect 7692 7588 7696 7644
rect 7696 7588 7752 7644
rect 7752 7588 7756 7644
rect 7692 7584 7756 7588
rect 7772 7644 7836 7648
rect 7772 7588 7776 7644
rect 7776 7588 7832 7644
rect 7832 7588 7836 7644
rect 7772 7584 7836 7588
rect 7852 7644 7916 7648
rect 7852 7588 7856 7644
rect 7856 7588 7912 7644
rect 7912 7588 7916 7644
rect 7852 7584 7916 7588
rect 5948 7516 6012 7580
rect 12612 7644 12676 7648
rect 12612 7588 12616 7644
rect 12616 7588 12672 7644
rect 12672 7588 12676 7644
rect 12612 7584 12676 7588
rect 12692 7644 12756 7648
rect 12692 7588 12696 7644
rect 12696 7588 12752 7644
rect 12752 7588 12756 7644
rect 12692 7584 12756 7588
rect 12772 7644 12836 7648
rect 12772 7588 12776 7644
rect 12776 7588 12832 7644
rect 12832 7588 12836 7644
rect 12772 7584 12836 7588
rect 12852 7644 12916 7648
rect 12852 7588 12856 7644
rect 12856 7588 12912 7644
rect 12912 7588 12916 7644
rect 12852 7584 12916 7588
rect 17612 7644 17676 7648
rect 17612 7588 17616 7644
rect 17616 7588 17672 7644
rect 17672 7588 17676 7644
rect 17612 7584 17676 7588
rect 17692 7644 17756 7648
rect 17692 7588 17696 7644
rect 17696 7588 17752 7644
rect 17752 7588 17756 7644
rect 17692 7584 17756 7588
rect 17772 7644 17836 7648
rect 17772 7588 17776 7644
rect 17776 7588 17832 7644
rect 17832 7588 17836 7644
rect 17772 7584 17836 7588
rect 17852 7644 17916 7648
rect 17852 7588 17856 7644
rect 17856 7588 17912 7644
rect 17912 7588 17916 7644
rect 17852 7584 17916 7588
rect 5028 7380 5092 7444
rect 8340 7380 8404 7444
rect 3556 7244 3620 7308
rect 6132 7244 6196 7308
rect 10732 7244 10796 7308
rect 1716 7168 1780 7172
rect 1716 7112 1766 7168
rect 1766 7112 1780 7168
rect 1716 7108 1780 7112
rect 10364 7108 10428 7172
rect 12388 7108 12452 7172
rect 1952 7100 2016 7104
rect 1952 7044 1956 7100
rect 1956 7044 2012 7100
rect 2012 7044 2016 7100
rect 1952 7040 2016 7044
rect 2032 7100 2096 7104
rect 2032 7044 2036 7100
rect 2036 7044 2092 7100
rect 2092 7044 2096 7100
rect 2032 7040 2096 7044
rect 2112 7100 2176 7104
rect 2112 7044 2116 7100
rect 2116 7044 2172 7100
rect 2172 7044 2176 7100
rect 2112 7040 2176 7044
rect 2192 7100 2256 7104
rect 2192 7044 2196 7100
rect 2196 7044 2252 7100
rect 2252 7044 2256 7100
rect 2192 7040 2256 7044
rect 6952 7100 7016 7104
rect 6952 7044 6956 7100
rect 6956 7044 7012 7100
rect 7012 7044 7016 7100
rect 6952 7040 7016 7044
rect 7032 7100 7096 7104
rect 7032 7044 7036 7100
rect 7036 7044 7092 7100
rect 7092 7044 7096 7100
rect 7032 7040 7096 7044
rect 7112 7100 7176 7104
rect 7112 7044 7116 7100
rect 7116 7044 7172 7100
rect 7172 7044 7176 7100
rect 7112 7040 7176 7044
rect 7192 7100 7256 7104
rect 7192 7044 7196 7100
rect 7196 7044 7252 7100
rect 7252 7044 7256 7100
rect 7192 7040 7256 7044
rect 11952 7100 12016 7104
rect 11952 7044 11956 7100
rect 11956 7044 12012 7100
rect 12012 7044 12016 7100
rect 11952 7040 12016 7044
rect 12032 7100 12096 7104
rect 12032 7044 12036 7100
rect 12036 7044 12092 7100
rect 12092 7044 12096 7100
rect 12032 7040 12096 7044
rect 12112 7100 12176 7104
rect 12112 7044 12116 7100
rect 12116 7044 12172 7100
rect 12172 7044 12176 7100
rect 12112 7040 12176 7044
rect 12192 7100 12256 7104
rect 12192 7044 12196 7100
rect 12196 7044 12252 7100
rect 12252 7044 12256 7100
rect 12192 7040 12256 7044
rect 16952 7100 17016 7104
rect 16952 7044 16956 7100
rect 16956 7044 17012 7100
rect 17012 7044 17016 7100
rect 16952 7040 17016 7044
rect 17032 7100 17096 7104
rect 17032 7044 17036 7100
rect 17036 7044 17092 7100
rect 17092 7044 17096 7100
rect 17032 7040 17096 7044
rect 17112 7100 17176 7104
rect 17112 7044 17116 7100
rect 17116 7044 17172 7100
rect 17172 7044 17176 7100
rect 17112 7040 17176 7044
rect 17192 7100 17256 7104
rect 17192 7044 17196 7100
rect 17196 7044 17252 7100
rect 17252 7044 17256 7100
rect 17192 7040 17256 7044
rect 3924 7032 3988 7036
rect 3924 6976 3938 7032
rect 3938 6976 3988 7032
rect 3924 6972 3988 6976
rect 9444 6972 9508 7036
rect 11100 7032 11164 7036
rect 11100 6976 11114 7032
rect 11114 6976 11164 7032
rect 11100 6972 11164 6976
rect 3372 6836 3436 6900
rect 13124 6836 13188 6900
rect 6500 6700 6564 6764
rect 15700 6700 15764 6764
rect 2612 6556 2676 6560
rect 2612 6500 2616 6556
rect 2616 6500 2672 6556
rect 2672 6500 2676 6556
rect 2612 6496 2676 6500
rect 2692 6556 2756 6560
rect 2692 6500 2696 6556
rect 2696 6500 2752 6556
rect 2752 6500 2756 6556
rect 2692 6496 2756 6500
rect 2772 6556 2836 6560
rect 2772 6500 2776 6556
rect 2776 6500 2832 6556
rect 2832 6500 2836 6556
rect 2772 6496 2836 6500
rect 2852 6556 2916 6560
rect 2852 6500 2856 6556
rect 2856 6500 2912 6556
rect 2912 6500 2916 6556
rect 2852 6496 2916 6500
rect 7612 6556 7676 6560
rect 7612 6500 7616 6556
rect 7616 6500 7672 6556
rect 7672 6500 7676 6556
rect 7612 6496 7676 6500
rect 7692 6556 7756 6560
rect 7692 6500 7696 6556
rect 7696 6500 7752 6556
rect 7752 6500 7756 6556
rect 7692 6496 7756 6500
rect 7772 6556 7836 6560
rect 7772 6500 7776 6556
rect 7776 6500 7832 6556
rect 7832 6500 7836 6556
rect 7772 6496 7836 6500
rect 7852 6556 7916 6560
rect 7852 6500 7856 6556
rect 7856 6500 7912 6556
rect 7912 6500 7916 6556
rect 7852 6496 7916 6500
rect 12612 6556 12676 6560
rect 12612 6500 12616 6556
rect 12616 6500 12672 6556
rect 12672 6500 12676 6556
rect 12612 6496 12676 6500
rect 12692 6556 12756 6560
rect 12692 6500 12696 6556
rect 12696 6500 12752 6556
rect 12752 6500 12756 6556
rect 12692 6496 12756 6500
rect 12772 6556 12836 6560
rect 12772 6500 12776 6556
rect 12776 6500 12832 6556
rect 12832 6500 12836 6556
rect 12772 6496 12836 6500
rect 12852 6556 12916 6560
rect 12852 6500 12856 6556
rect 12856 6500 12912 6556
rect 12912 6500 12916 6556
rect 12852 6496 12916 6500
rect 17612 6556 17676 6560
rect 17612 6500 17616 6556
rect 17616 6500 17672 6556
rect 17672 6500 17676 6556
rect 17612 6496 17676 6500
rect 17692 6556 17756 6560
rect 17692 6500 17696 6556
rect 17696 6500 17752 6556
rect 17752 6500 17756 6556
rect 17692 6496 17756 6500
rect 17772 6556 17836 6560
rect 17772 6500 17776 6556
rect 17776 6500 17832 6556
rect 17832 6500 17836 6556
rect 17772 6496 17836 6500
rect 17852 6556 17916 6560
rect 17852 6500 17856 6556
rect 17856 6500 17912 6556
rect 17912 6500 17916 6556
rect 17852 6496 17916 6500
rect 1532 6428 1596 6492
rect 10180 6428 10244 6492
rect 13676 6428 13740 6492
rect 15700 6428 15764 6492
rect 8156 6292 8220 6356
rect 10364 6292 10428 6356
rect 4292 6156 4356 6220
rect 4660 6156 4724 6220
rect 6500 6156 6564 6220
rect 1952 6012 2016 6016
rect 1952 5956 1956 6012
rect 1956 5956 2012 6012
rect 2012 5956 2016 6012
rect 1952 5952 2016 5956
rect 2032 6012 2096 6016
rect 2032 5956 2036 6012
rect 2036 5956 2092 6012
rect 2092 5956 2096 6012
rect 2032 5952 2096 5956
rect 2112 6012 2176 6016
rect 2112 5956 2116 6012
rect 2116 5956 2172 6012
rect 2172 5956 2176 6012
rect 2112 5952 2176 5956
rect 2192 6012 2256 6016
rect 2192 5956 2196 6012
rect 2196 5956 2252 6012
rect 2252 5956 2256 6012
rect 2192 5952 2256 5956
rect 4108 5944 4172 5948
rect 4108 5888 4122 5944
rect 4122 5888 4172 5944
rect 4108 5884 4172 5888
rect 5948 5884 6012 5948
rect 4844 5748 4908 5812
rect 5764 5748 5828 5812
rect 11468 6020 11532 6084
rect 6952 6012 7016 6016
rect 6952 5956 6956 6012
rect 6956 5956 7012 6012
rect 7012 5956 7016 6012
rect 6952 5952 7016 5956
rect 7032 6012 7096 6016
rect 7032 5956 7036 6012
rect 7036 5956 7092 6012
rect 7092 5956 7096 6012
rect 7032 5952 7096 5956
rect 7112 6012 7176 6016
rect 7112 5956 7116 6012
rect 7116 5956 7172 6012
rect 7172 5956 7176 6012
rect 7112 5952 7176 5956
rect 7192 6012 7256 6016
rect 7192 5956 7196 6012
rect 7196 5956 7252 6012
rect 7252 5956 7256 6012
rect 7192 5952 7256 5956
rect 11952 6012 12016 6016
rect 11952 5956 11956 6012
rect 11956 5956 12012 6012
rect 12012 5956 12016 6012
rect 11952 5952 12016 5956
rect 12032 6012 12096 6016
rect 12032 5956 12036 6012
rect 12036 5956 12092 6012
rect 12092 5956 12096 6012
rect 12032 5952 12096 5956
rect 12112 6012 12176 6016
rect 12112 5956 12116 6012
rect 12116 5956 12172 6012
rect 12172 5956 12176 6012
rect 12112 5952 12176 5956
rect 12192 6012 12256 6016
rect 12192 5956 12196 6012
rect 12196 5956 12252 6012
rect 12252 5956 12256 6012
rect 12192 5952 12256 5956
rect 16952 6012 17016 6016
rect 16952 5956 16956 6012
rect 16956 5956 17012 6012
rect 17012 5956 17016 6012
rect 16952 5952 17016 5956
rect 17032 6012 17096 6016
rect 17032 5956 17036 6012
rect 17036 5956 17092 6012
rect 17092 5956 17096 6012
rect 17032 5952 17096 5956
rect 17112 6012 17176 6016
rect 17112 5956 17116 6012
rect 17116 5956 17172 6012
rect 17172 5956 17176 6012
rect 17112 5952 17176 5956
rect 17192 6012 17256 6016
rect 17192 5956 17196 6012
rect 17196 5956 17252 6012
rect 17252 5956 17256 6012
rect 17192 5952 17256 5956
rect 8156 5884 8220 5948
rect 9812 5884 9876 5948
rect 10732 5748 10796 5812
rect 18092 5748 18156 5812
rect 796 5612 860 5676
rect 9996 5476 10060 5540
rect 11284 5476 11348 5540
rect 18276 5612 18340 5676
rect 18460 5476 18524 5540
rect 2612 5468 2676 5472
rect 2612 5412 2616 5468
rect 2616 5412 2672 5468
rect 2672 5412 2676 5468
rect 2612 5408 2676 5412
rect 2692 5468 2756 5472
rect 2692 5412 2696 5468
rect 2696 5412 2752 5468
rect 2752 5412 2756 5468
rect 2692 5408 2756 5412
rect 2772 5468 2836 5472
rect 2772 5412 2776 5468
rect 2776 5412 2832 5468
rect 2832 5412 2836 5468
rect 2772 5408 2836 5412
rect 2852 5468 2916 5472
rect 2852 5412 2856 5468
rect 2856 5412 2912 5468
rect 2912 5412 2916 5468
rect 2852 5408 2916 5412
rect 7612 5468 7676 5472
rect 7612 5412 7616 5468
rect 7616 5412 7672 5468
rect 7672 5412 7676 5468
rect 7612 5408 7676 5412
rect 7692 5468 7756 5472
rect 7692 5412 7696 5468
rect 7696 5412 7752 5468
rect 7752 5412 7756 5468
rect 7692 5408 7756 5412
rect 7772 5468 7836 5472
rect 7772 5412 7776 5468
rect 7776 5412 7832 5468
rect 7832 5412 7836 5468
rect 7772 5408 7836 5412
rect 7852 5468 7916 5472
rect 7852 5412 7856 5468
rect 7856 5412 7912 5468
rect 7912 5412 7916 5468
rect 7852 5408 7916 5412
rect 12612 5468 12676 5472
rect 12612 5412 12616 5468
rect 12616 5412 12672 5468
rect 12672 5412 12676 5468
rect 12612 5408 12676 5412
rect 12692 5468 12756 5472
rect 12692 5412 12696 5468
rect 12696 5412 12752 5468
rect 12752 5412 12756 5468
rect 12692 5408 12756 5412
rect 12772 5468 12836 5472
rect 12772 5412 12776 5468
rect 12776 5412 12832 5468
rect 12832 5412 12836 5468
rect 12772 5408 12836 5412
rect 12852 5468 12916 5472
rect 12852 5412 12856 5468
rect 12856 5412 12912 5468
rect 12912 5412 12916 5468
rect 12852 5408 12916 5412
rect 17612 5468 17676 5472
rect 17612 5412 17616 5468
rect 17616 5412 17672 5468
rect 17672 5412 17676 5468
rect 17612 5408 17676 5412
rect 17692 5468 17756 5472
rect 17692 5412 17696 5468
rect 17696 5412 17752 5468
rect 17752 5412 17756 5468
rect 17692 5408 17756 5412
rect 17772 5468 17836 5472
rect 17772 5412 17776 5468
rect 17776 5412 17832 5468
rect 17832 5412 17836 5468
rect 17772 5408 17836 5412
rect 17852 5468 17916 5472
rect 17852 5412 17856 5468
rect 17856 5412 17912 5468
rect 17912 5412 17916 5468
rect 17852 5408 17916 5412
rect 11284 5340 11348 5404
rect 12388 5340 12452 5404
rect 3004 5264 3068 5268
rect 3004 5208 3054 5264
rect 3054 5208 3068 5264
rect 3004 5204 3068 5208
rect 5580 5204 5644 5268
rect 6684 5204 6748 5268
rect 9076 5204 9140 5268
rect 980 5068 1044 5132
rect 9628 5068 9692 5132
rect 13308 5204 13372 5268
rect 6316 4932 6380 4996
rect 7420 4932 7484 4996
rect 1952 4924 2016 4928
rect 1952 4868 1956 4924
rect 1956 4868 2012 4924
rect 2012 4868 2016 4924
rect 1952 4864 2016 4868
rect 2032 4924 2096 4928
rect 2032 4868 2036 4924
rect 2036 4868 2092 4924
rect 2092 4868 2096 4924
rect 2032 4864 2096 4868
rect 2112 4924 2176 4928
rect 2112 4868 2116 4924
rect 2116 4868 2172 4924
rect 2172 4868 2176 4924
rect 2112 4864 2176 4868
rect 2192 4924 2256 4928
rect 2192 4868 2196 4924
rect 2196 4868 2252 4924
rect 2252 4868 2256 4924
rect 2192 4864 2256 4868
rect 6952 4924 7016 4928
rect 6952 4868 6956 4924
rect 6956 4868 7012 4924
rect 7012 4868 7016 4924
rect 6952 4864 7016 4868
rect 7032 4924 7096 4928
rect 7032 4868 7036 4924
rect 7036 4868 7092 4924
rect 7092 4868 7096 4924
rect 7032 4864 7096 4868
rect 7112 4924 7176 4928
rect 7112 4868 7116 4924
rect 7116 4868 7172 4924
rect 7172 4868 7176 4924
rect 7112 4864 7176 4868
rect 7192 4924 7256 4928
rect 7192 4868 7196 4924
rect 7196 4868 7252 4924
rect 7252 4868 7256 4924
rect 7192 4864 7256 4868
rect 11952 4924 12016 4928
rect 11952 4868 11956 4924
rect 11956 4868 12012 4924
rect 12012 4868 12016 4924
rect 11952 4864 12016 4868
rect 12032 4924 12096 4928
rect 12032 4868 12036 4924
rect 12036 4868 12092 4924
rect 12092 4868 12096 4924
rect 12032 4864 12096 4868
rect 12112 4924 12176 4928
rect 12112 4868 12116 4924
rect 12116 4868 12172 4924
rect 12172 4868 12176 4924
rect 12112 4864 12176 4868
rect 12192 4924 12256 4928
rect 12192 4868 12196 4924
rect 12196 4868 12252 4924
rect 12252 4868 12256 4924
rect 12192 4864 12256 4868
rect 16952 4924 17016 4928
rect 16952 4868 16956 4924
rect 16956 4868 17012 4924
rect 17012 4868 17016 4924
rect 16952 4864 17016 4868
rect 17032 4924 17096 4928
rect 17032 4868 17036 4924
rect 17036 4868 17092 4924
rect 17092 4868 17096 4924
rect 17032 4864 17096 4868
rect 17112 4924 17176 4928
rect 17112 4868 17116 4924
rect 17116 4868 17172 4924
rect 17172 4868 17176 4924
rect 17112 4864 17176 4868
rect 17192 4924 17256 4928
rect 17192 4868 17196 4924
rect 17196 4868 17252 4924
rect 17252 4868 17256 4924
rect 17192 4864 17256 4868
rect 5212 4796 5276 4860
rect 14780 4856 14844 4860
rect 14780 4800 14830 4856
rect 14830 4800 14844 4856
rect 14780 4796 14844 4800
rect 5028 4524 5092 4588
rect 15148 4660 15212 4724
rect 16436 4524 16500 4588
rect 6132 4388 6196 4452
rect 7420 4388 7484 4452
rect 13492 4448 13556 4452
rect 13492 4392 13542 4448
rect 13542 4392 13556 4448
rect 13492 4388 13556 4392
rect 13676 4388 13740 4452
rect 2612 4380 2676 4384
rect 2612 4324 2616 4380
rect 2616 4324 2672 4380
rect 2672 4324 2676 4380
rect 2612 4320 2676 4324
rect 2692 4380 2756 4384
rect 2692 4324 2696 4380
rect 2696 4324 2752 4380
rect 2752 4324 2756 4380
rect 2692 4320 2756 4324
rect 2772 4380 2836 4384
rect 2772 4324 2776 4380
rect 2776 4324 2832 4380
rect 2832 4324 2836 4380
rect 2772 4320 2836 4324
rect 2852 4380 2916 4384
rect 2852 4324 2856 4380
rect 2856 4324 2912 4380
rect 2912 4324 2916 4380
rect 2852 4320 2916 4324
rect 7612 4380 7676 4384
rect 7612 4324 7616 4380
rect 7616 4324 7672 4380
rect 7672 4324 7676 4380
rect 7612 4320 7676 4324
rect 7692 4380 7756 4384
rect 7692 4324 7696 4380
rect 7696 4324 7752 4380
rect 7752 4324 7756 4380
rect 7692 4320 7756 4324
rect 7772 4380 7836 4384
rect 7772 4324 7776 4380
rect 7776 4324 7832 4380
rect 7832 4324 7836 4380
rect 7772 4320 7836 4324
rect 7852 4380 7916 4384
rect 7852 4324 7856 4380
rect 7856 4324 7912 4380
rect 7912 4324 7916 4380
rect 7852 4320 7916 4324
rect 12612 4380 12676 4384
rect 12612 4324 12616 4380
rect 12616 4324 12672 4380
rect 12672 4324 12676 4380
rect 12612 4320 12676 4324
rect 12692 4380 12756 4384
rect 12692 4324 12696 4380
rect 12696 4324 12752 4380
rect 12752 4324 12756 4380
rect 12692 4320 12756 4324
rect 12772 4380 12836 4384
rect 12772 4324 12776 4380
rect 12776 4324 12832 4380
rect 12832 4324 12836 4380
rect 12772 4320 12836 4324
rect 12852 4380 12916 4384
rect 12852 4324 12856 4380
rect 12856 4324 12912 4380
rect 12912 4324 12916 4380
rect 12852 4320 12916 4324
rect 17612 4380 17676 4384
rect 17612 4324 17616 4380
rect 17616 4324 17672 4380
rect 17672 4324 17676 4380
rect 17612 4320 17676 4324
rect 17692 4380 17756 4384
rect 17692 4324 17696 4380
rect 17696 4324 17752 4380
rect 17752 4324 17756 4380
rect 17692 4320 17756 4324
rect 17772 4380 17836 4384
rect 17772 4324 17776 4380
rect 17776 4324 17832 4380
rect 17832 4324 17836 4380
rect 17772 4320 17836 4324
rect 17852 4380 17916 4384
rect 17852 4324 17856 4380
rect 17856 4324 17912 4380
rect 17912 4324 17916 4380
rect 17852 4320 17916 4324
rect 3188 4252 3252 4316
rect 8340 4116 8404 4180
rect 11100 4252 11164 4316
rect 10732 3980 10796 4044
rect 11652 3980 11716 4044
rect 14964 4116 15028 4180
rect 15148 4116 15212 4180
rect 16068 4176 16132 4180
rect 16068 4120 16082 4176
rect 16082 4120 16132 4176
rect 16068 4116 16132 4120
rect 14044 3980 14108 4044
rect 18828 3980 18892 4044
rect 4476 3844 4540 3908
rect 6316 3844 6380 3908
rect 8524 3904 8588 3908
rect 8524 3848 8574 3904
rect 8574 3848 8588 3904
rect 8524 3844 8588 3848
rect 1952 3836 2016 3840
rect 1952 3780 1956 3836
rect 1956 3780 2012 3836
rect 2012 3780 2016 3836
rect 1952 3776 2016 3780
rect 2032 3836 2096 3840
rect 2032 3780 2036 3836
rect 2036 3780 2092 3836
rect 2092 3780 2096 3836
rect 2032 3776 2096 3780
rect 2112 3836 2176 3840
rect 2112 3780 2116 3836
rect 2116 3780 2172 3836
rect 2172 3780 2176 3836
rect 2112 3776 2176 3780
rect 2192 3836 2256 3840
rect 2192 3780 2196 3836
rect 2196 3780 2252 3836
rect 2252 3780 2256 3836
rect 2192 3776 2256 3780
rect 6952 3836 7016 3840
rect 6952 3780 6956 3836
rect 6956 3780 7012 3836
rect 7012 3780 7016 3836
rect 6952 3776 7016 3780
rect 7032 3836 7096 3840
rect 7032 3780 7036 3836
rect 7036 3780 7092 3836
rect 7092 3780 7096 3836
rect 7032 3776 7096 3780
rect 7112 3836 7176 3840
rect 7112 3780 7116 3836
rect 7116 3780 7172 3836
rect 7172 3780 7176 3836
rect 7112 3776 7176 3780
rect 7192 3836 7256 3840
rect 7192 3780 7196 3836
rect 7196 3780 7252 3836
rect 7252 3780 7256 3836
rect 7192 3776 7256 3780
rect 11952 3836 12016 3840
rect 11952 3780 11956 3836
rect 11956 3780 12012 3836
rect 12012 3780 12016 3836
rect 11952 3776 12016 3780
rect 12032 3836 12096 3840
rect 12032 3780 12036 3836
rect 12036 3780 12092 3836
rect 12092 3780 12096 3836
rect 12032 3776 12096 3780
rect 12112 3836 12176 3840
rect 12112 3780 12116 3836
rect 12116 3780 12172 3836
rect 12172 3780 12176 3836
rect 12112 3776 12176 3780
rect 12192 3836 12256 3840
rect 12192 3780 12196 3836
rect 12196 3780 12252 3836
rect 12252 3780 12256 3836
rect 12192 3776 12256 3780
rect 16952 3836 17016 3840
rect 16952 3780 16956 3836
rect 16956 3780 17012 3836
rect 17012 3780 17016 3836
rect 16952 3776 17016 3780
rect 17032 3836 17096 3840
rect 17032 3780 17036 3836
rect 17036 3780 17092 3836
rect 17092 3780 17096 3836
rect 17032 3776 17096 3780
rect 17112 3836 17176 3840
rect 17112 3780 17116 3836
rect 17116 3780 17172 3836
rect 17172 3780 17176 3836
rect 17112 3776 17176 3780
rect 17192 3836 17256 3840
rect 17192 3780 17196 3836
rect 17196 3780 17252 3836
rect 17252 3780 17256 3836
rect 17192 3776 17256 3780
rect 3372 3436 3436 3500
rect 4108 3436 4172 3500
rect 5948 3572 6012 3636
rect 9260 3708 9324 3772
rect 13860 3572 13924 3636
rect 6500 3300 6564 3364
rect 9260 3300 9324 3364
rect 16804 3360 16868 3364
rect 16804 3304 16854 3360
rect 16854 3304 16868 3360
rect 16804 3300 16868 3304
rect 2612 3292 2676 3296
rect 2612 3236 2616 3292
rect 2616 3236 2672 3292
rect 2672 3236 2676 3292
rect 2612 3232 2676 3236
rect 2692 3292 2756 3296
rect 2692 3236 2696 3292
rect 2696 3236 2752 3292
rect 2752 3236 2756 3292
rect 2692 3232 2756 3236
rect 2772 3292 2836 3296
rect 2772 3236 2776 3292
rect 2776 3236 2832 3292
rect 2832 3236 2836 3292
rect 2772 3232 2836 3236
rect 2852 3292 2916 3296
rect 2852 3236 2856 3292
rect 2856 3236 2912 3292
rect 2912 3236 2916 3292
rect 2852 3232 2916 3236
rect 7612 3292 7676 3296
rect 7612 3236 7616 3292
rect 7616 3236 7672 3292
rect 7672 3236 7676 3292
rect 7612 3232 7676 3236
rect 7692 3292 7756 3296
rect 7692 3236 7696 3292
rect 7696 3236 7752 3292
rect 7752 3236 7756 3292
rect 7692 3232 7756 3236
rect 7772 3292 7836 3296
rect 7772 3236 7776 3292
rect 7776 3236 7832 3292
rect 7832 3236 7836 3292
rect 7772 3232 7836 3236
rect 7852 3292 7916 3296
rect 7852 3236 7856 3292
rect 7856 3236 7912 3292
rect 7912 3236 7916 3292
rect 7852 3232 7916 3236
rect 12612 3292 12676 3296
rect 12612 3236 12616 3292
rect 12616 3236 12672 3292
rect 12672 3236 12676 3292
rect 12612 3232 12676 3236
rect 12692 3292 12756 3296
rect 12692 3236 12696 3292
rect 12696 3236 12752 3292
rect 12752 3236 12756 3292
rect 12692 3232 12756 3236
rect 12772 3292 12836 3296
rect 12772 3236 12776 3292
rect 12776 3236 12832 3292
rect 12832 3236 12836 3292
rect 12772 3232 12836 3236
rect 12852 3292 12916 3296
rect 12852 3236 12856 3292
rect 12856 3236 12912 3292
rect 12912 3236 12916 3292
rect 12852 3232 12916 3236
rect 17612 3292 17676 3296
rect 17612 3236 17616 3292
rect 17616 3236 17672 3292
rect 17672 3236 17676 3292
rect 17612 3232 17676 3236
rect 17692 3292 17756 3296
rect 17692 3236 17696 3292
rect 17696 3236 17752 3292
rect 17752 3236 17756 3292
rect 17692 3232 17756 3236
rect 17772 3292 17836 3296
rect 17772 3236 17776 3292
rect 17776 3236 17832 3292
rect 17832 3236 17836 3292
rect 17772 3232 17836 3236
rect 17852 3292 17916 3296
rect 17852 3236 17856 3292
rect 17856 3236 17912 3292
rect 17912 3236 17916 3292
rect 17852 3232 17916 3236
rect 11284 3164 11348 3228
rect 3740 3028 3804 3092
rect 2452 2892 2516 2956
rect 1952 2748 2016 2752
rect 1952 2692 1956 2748
rect 1956 2692 2012 2748
rect 2012 2692 2016 2748
rect 1952 2688 2016 2692
rect 2032 2748 2096 2752
rect 2032 2692 2036 2748
rect 2036 2692 2092 2748
rect 2092 2692 2096 2748
rect 2032 2688 2096 2692
rect 2112 2748 2176 2752
rect 2112 2692 2116 2748
rect 2116 2692 2172 2748
rect 2172 2692 2176 2748
rect 2112 2688 2176 2692
rect 2192 2748 2256 2752
rect 2192 2692 2196 2748
rect 2196 2692 2252 2748
rect 2252 2692 2256 2748
rect 2192 2688 2256 2692
rect 6952 2748 7016 2752
rect 6952 2692 6956 2748
rect 6956 2692 7012 2748
rect 7012 2692 7016 2748
rect 6952 2688 7016 2692
rect 7032 2748 7096 2752
rect 7032 2692 7036 2748
rect 7036 2692 7092 2748
rect 7092 2692 7096 2748
rect 7032 2688 7096 2692
rect 7112 2748 7176 2752
rect 7112 2692 7116 2748
rect 7116 2692 7172 2748
rect 7172 2692 7176 2748
rect 7112 2688 7176 2692
rect 7192 2748 7256 2752
rect 7192 2692 7196 2748
rect 7196 2692 7252 2748
rect 7252 2692 7256 2748
rect 7192 2688 7256 2692
rect 3556 2620 3620 2684
rect 1348 2484 1412 2548
rect 11952 2748 12016 2752
rect 11952 2692 11956 2748
rect 11956 2692 12012 2748
rect 12012 2692 12016 2748
rect 11952 2688 12016 2692
rect 12032 2748 12096 2752
rect 12032 2692 12036 2748
rect 12036 2692 12092 2748
rect 12092 2692 12096 2748
rect 12032 2688 12096 2692
rect 12112 2748 12176 2752
rect 12112 2692 12116 2748
rect 12116 2692 12172 2748
rect 12172 2692 12176 2748
rect 12112 2688 12176 2692
rect 12192 2748 12256 2752
rect 12192 2692 12196 2748
rect 12196 2692 12252 2748
rect 12252 2692 12256 2748
rect 12192 2688 12256 2692
rect 16952 2748 17016 2752
rect 16952 2692 16956 2748
rect 16956 2692 17012 2748
rect 17012 2692 17016 2748
rect 16952 2688 17016 2692
rect 17032 2748 17096 2752
rect 17032 2692 17036 2748
rect 17036 2692 17092 2748
rect 17092 2692 17096 2748
rect 17032 2688 17096 2692
rect 17112 2748 17176 2752
rect 17112 2692 17116 2748
rect 17116 2692 17172 2748
rect 17172 2692 17176 2748
rect 17112 2688 17176 2692
rect 17192 2748 17256 2752
rect 17192 2692 17196 2748
rect 17196 2692 17252 2748
rect 17252 2692 17256 2748
rect 17192 2688 17256 2692
rect 8156 2680 8220 2684
rect 8156 2624 8206 2680
rect 8206 2624 8220 2680
rect 8156 2620 8220 2624
rect 8708 2680 8772 2684
rect 8708 2624 8722 2680
rect 8722 2624 8772 2680
rect 8708 2620 8772 2624
rect 8892 2620 8956 2684
rect 16252 2620 16316 2684
rect 10364 2484 10428 2548
rect 10916 2484 10980 2548
rect 16620 2484 16684 2548
rect 14412 2348 14476 2412
rect 18644 2348 18708 2412
rect 5396 2212 5460 2276
rect 2612 2204 2676 2208
rect 2612 2148 2616 2204
rect 2616 2148 2672 2204
rect 2672 2148 2676 2204
rect 2612 2144 2676 2148
rect 2692 2204 2756 2208
rect 2692 2148 2696 2204
rect 2696 2148 2752 2204
rect 2752 2148 2756 2204
rect 2692 2144 2756 2148
rect 2772 2204 2836 2208
rect 2772 2148 2776 2204
rect 2776 2148 2832 2204
rect 2832 2148 2836 2204
rect 2772 2144 2836 2148
rect 2852 2204 2916 2208
rect 2852 2148 2856 2204
rect 2856 2148 2912 2204
rect 2912 2148 2916 2204
rect 2852 2144 2916 2148
rect 7612 2204 7676 2208
rect 7612 2148 7616 2204
rect 7616 2148 7672 2204
rect 7672 2148 7676 2204
rect 7612 2144 7676 2148
rect 7692 2204 7756 2208
rect 7692 2148 7696 2204
rect 7696 2148 7752 2204
rect 7752 2148 7756 2204
rect 7692 2144 7756 2148
rect 7772 2204 7836 2208
rect 7772 2148 7776 2204
rect 7776 2148 7832 2204
rect 7832 2148 7836 2204
rect 7772 2144 7836 2148
rect 7852 2204 7916 2208
rect 7852 2148 7856 2204
rect 7856 2148 7912 2204
rect 7912 2148 7916 2204
rect 7852 2144 7916 2148
rect 12612 2204 12676 2208
rect 12612 2148 12616 2204
rect 12616 2148 12672 2204
rect 12672 2148 12676 2204
rect 12612 2144 12676 2148
rect 12692 2204 12756 2208
rect 12692 2148 12696 2204
rect 12696 2148 12752 2204
rect 12752 2148 12756 2204
rect 12692 2144 12756 2148
rect 12772 2204 12836 2208
rect 12772 2148 12776 2204
rect 12776 2148 12832 2204
rect 12832 2148 12836 2204
rect 12772 2144 12836 2148
rect 12852 2204 12916 2208
rect 12852 2148 12856 2204
rect 12856 2148 12912 2204
rect 12912 2148 12916 2204
rect 12852 2144 12916 2148
rect 17612 2204 17676 2208
rect 17612 2148 17616 2204
rect 17616 2148 17672 2204
rect 17672 2148 17676 2204
rect 17612 2144 17676 2148
rect 17692 2204 17756 2208
rect 17692 2148 17696 2204
rect 17696 2148 17752 2204
rect 17752 2148 17756 2204
rect 17692 2144 17756 2148
rect 17772 2204 17836 2208
rect 17772 2148 17776 2204
rect 17776 2148 17832 2204
rect 17832 2148 17836 2204
rect 17772 2144 17836 2148
rect 17852 2204 17916 2208
rect 17852 2148 17856 2204
rect 17856 2148 17912 2204
rect 17912 2148 17916 2204
rect 17852 2144 17916 2148
rect 10548 1804 10612 1868
rect 15332 1940 15396 2004
rect 17908 1668 17972 1732
rect 19012 1668 19076 1732
rect 17908 1396 17972 1460
rect 1716 988 1780 1052
rect 3924 852 3988 916
rect 796 716 860 780
rect 4660 580 4724 644
rect 13124 444 13188 508
<< metal4 >>
rect 15883 18732 15949 18733
rect 15883 18668 15884 18732
rect 15948 18668 15949 18732
rect 15883 18667 15949 18668
rect 5027 18596 5093 18597
rect 5027 18532 5028 18596
rect 5092 18532 5093 18596
rect 5027 18531 5093 18532
rect 1531 18460 1597 18461
rect 1531 18396 1532 18460
rect 1596 18396 1597 18460
rect 1531 18395 1597 18396
rect 795 15332 861 15333
rect 795 15268 796 15332
rect 860 15268 861 15332
rect 795 15267 861 15268
rect 798 9077 858 15267
rect 795 9076 861 9077
rect 795 9012 796 9076
rect 860 9012 861 9076
rect 795 9011 861 9012
rect 798 5677 858 9011
rect 795 5676 861 5677
rect 795 5612 796 5676
rect 860 5612 861 5676
rect 795 5611 861 5612
rect 982 5133 1042 16542
rect 1163 13836 1229 13837
rect 1163 13772 1164 13836
rect 1228 13772 1229 13836
rect 1163 13771 1229 13772
rect 979 5132 1045 5133
rect 979 5068 980 5132
rect 1044 5068 1045 5132
rect 979 5067 1045 5068
rect 1166 2790 1226 13771
rect 1347 13428 1413 13429
rect 1347 13364 1348 13428
rect 1412 13364 1413 13428
rect 1347 13363 1413 13364
rect 1350 8533 1410 13363
rect 1534 8669 1594 18395
rect 1944 16896 2264 17456
rect 2604 17440 2924 17456
rect 2604 17376 2612 17440
rect 2676 17376 2692 17440
rect 2756 17376 2772 17440
rect 2836 17376 2852 17440
rect 2916 17376 2924 17440
rect 2451 16964 2517 16965
rect 2451 16900 2452 16964
rect 2516 16900 2517 16964
rect 2451 16899 2517 16900
rect 1944 16832 1952 16896
rect 2016 16832 2032 16896
rect 2096 16832 2112 16896
rect 2176 16832 2192 16896
rect 2256 16832 2264 16896
rect 1944 15808 2264 16832
rect 1944 15744 1952 15808
rect 2016 15744 2032 15808
rect 2096 15744 2112 15808
rect 2176 15744 2192 15808
rect 2256 15744 2264 15808
rect 1944 14720 2264 15744
rect 1944 14656 1952 14720
rect 2016 14656 2032 14720
rect 2096 14656 2112 14720
rect 2176 14656 2192 14720
rect 2256 14656 2264 14720
rect 1944 13632 2264 14656
rect 2454 14245 2514 16899
rect 2604 16352 2924 17376
rect 3371 17100 3437 17101
rect 3371 17036 3372 17100
rect 3436 17036 3437 17100
rect 3371 17035 3437 17036
rect 2604 16288 2612 16352
rect 2676 16288 2692 16352
rect 2756 16288 2772 16352
rect 2836 16288 2852 16352
rect 2916 16288 2924 16352
rect 2604 15264 2924 16288
rect 2604 15200 2612 15264
rect 2676 15200 2692 15264
rect 2756 15200 2772 15264
rect 2836 15200 2852 15264
rect 2916 15200 2924 15264
rect 2451 14244 2517 14245
rect 2451 14180 2452 14244
rect 2516 14180 2517 14244
rect 2451 14179 2517 14180
rect 1944 13568 1952 13632
rect 2016 13568 2032 13632
rect 2096 13568 2112 13632
rect 2176 13568 2192 13632
rect 2256 13568 2264 13632
rect 1944 13294 2264 13568
rect 1944 13058 1986 13294
rect 2222 13058 2264 13294
rect 1944 12544 2264 13058
rect 1944 12480 1952 12544
rect 2016 12480 2032 12544
rect 2096 12480 2112 12544
rect 2176 12480 2192 12544
rect 2256 12480 2264 12544
rect 1944 11456 2264 12480
rect 2454 11525 2514 14179
rect 2604 14176 2924 15200
rect 2604 14112 2612 14176
rect 2676 14112 2692 14176
rect 2756 14112 2772 14176
rect 2836 14112 2852 14176
rect 2916 14112 2924 14176
rect 2604 13954 2924 14112
rect 2604 13718 2646 13954
rect 2882 13718 2924 13954
rect 2604 13088 2924 13718
rect 3187 13700 3253 13701
rect 3187 13636 3188 13700
rect 3252 13636 3253 13700
rect 3187 13635 3253 13636
rect 3003 13428 3069 13429
rect 3003 13364 3004 13428
rect 3068 13364 3069 13428
rect 3003 13363 3069 13364
rect 2604 13024 2612 13088
rect 2676 13024 2692 13088
rect 2756 13024 2772 13088
rect 2836 13024 2852 13088
rect 2916 13024 2924 13088
rect 2604 12000 2924 13024
rect 2604 11936 2612 12000
rect 2676 11936 2692 12000
rect 2756 11936 2772 12000
rect 2836 11936 2852 12000
rect 2916 11936 2924 12000
rect 2451 11524 2517 11525
rect 2451 11460 2452 11524
rect 2516 11460 2517 11524
rect 2451 11459 2517 11460
rect 1944 11392 1952 11456
rect 2016 11392 2032 11456
rect 2096 11392 2112 11456
rect 2176 11392 2192 11456
rect 2256 11392 2264 11456
rect 1944 10368 2264 11392
rect 1944 10304 1952 10368
rect 2016 10304 2032 10368
rect 2096 10304 2112 10368
rect 2176 10304 2192 10368
rect 2256 10304 2264 10368
rect 1715 9484 1781 9485
rect 1715 9420 1716 9484
rect 1780 9420 1781 9484
rect 1715 9419 1781 9420
rect 1531 8668 1597 8669
rect 1531 8604 1532 8668
rect 1596 8604 1597 8668
rect 1531 8603 1597 8604
rect 1347 8532 1413 8533
rect 1347 8468 1348 8532
rect 1412 8468 1413 8532
rect 1347 8467 1413 8468
rect 798 2730 1226 2790
rect 798 781 858 2730
rect 1350 2549 1410 8467
rect 1718 7850 1778 9419
rect 1488 7790 1778 7850
rect 1944 9280 2264 10304
rect 2604 10912 2924 11936
rect 2604 10848 2612 10912
rect 2676 10848 2692 10912
rect 2756 10848 2772 10912
rect 2836 10848 2852 10912
rect 2916 10848 2924 10912
rect 2604 9824 2924 10848
rect 3006 9893 3066 13363
rect 3190 10981 3250 13635
rect 3187 10980 3253 10981
rect 3187 10916 3188 10980
rect 3252 10916 3253 10980
rect 3187 10915 3253 10916
rect 3187 10164 3253 10165
rect 3187 10100 3188 10164
rect 3252 10100 3253 10164
rect 3187 10099 3253 10100
rect 3003 9892 3069 9893
rect 3003 9828 3004 9892
rect 3068 9828 3069 9892
rect 3003 9827 3069 9828
rect 2604 9760 2612 9824
rect 2676 9760 2692 9824
rect 2756 9760 2772 9824
rect 2836 9760 2852 9824
rect 2916 9760 2924 9824
rect 2451 9484 2517 9485
rect 2451 9420 2452 9484
rect 2516 9420 2517 9484
rect 2451 9419 2517 9420
rect 1944 9216 1952 9280
rect 2016 9216 2032 9280
rect 2096 9216 2112 9280
rect 2176 9216 2192 9280
rect 2256 9216 2264 9280
rect 1944 8294 2264 9216
rect 1944 8192 1986 8294
rect 2222 8192 2264 8294
rect 1944 8128 1952 8192
rect 2256 8128 2264 8192
rect 1944 8058 1986 8128
rect 2222 8058 2264 8128
rect 1488 6898 1548 7790
rect 1944 7104 2264 8058
rect 1944 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2264 7104
rect 1488 6838 1594 6898
rect 1534 6493 1594 6838
rect 1531 6492 1597 6493
rect 1531 6428 1532 6492
rect 1596 6428 1597 6492
rect 1531 6427 1597 6428
rect 1944 6016 2264 7040
rect 1944 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2264 6016
rect 1944 4928 2264 5952
rect 1944 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2264 4928
rect 1944 3840 2264 4864
rect 1944 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2264 3840
rect 1944 3294 2264 3776
rect 1944 3058 1986 3294
rect 2222 3058 2264 3294
rect 1944 2752 2264 3058
rect 2454 2957 2514 9419
rect 2604 8954 2924 9760
rect 3190 9485 3250 10099
rect 3374 9621 3434 17035
rect 4291 16012 4357 16013
rect 4291 15948 4292 16012
rect 4356 15948 4357 16012
rect 4291 15947 4357 15948
rect 4107 15332 4173 15333
rect 4107 15268 4108 15332
rect 4172 15268 4173 15332
rect 4107 15267 4173 15268
rect 3739 14652 3805 14653
rect 3739 14588 3740 14652
rect 3804 14588 3805 14652
rect 3739 14587 3805 14588
rect 3555 10844 3621 10845
rect 3555 10780 3556 10844
rect 3620 10780 3621 10844
rect 3555 10779 3621 10780
rect 3558 10437 3618 10779
rect 3742 10437 3802 14587
rect 3923 14244 3989 14245
rect 3923 14180 3924 14244
rect 3988 14180 3989 14244
rect 3923 14179 3989 14180
rect 3555 10436 3621 10437
rect 3555 10372 3556 10436
rect 3620 10372 3621 10436
rect 3555 10371 3621 10372
rect 3739 10436 3805 10437
rect 3739 10372 3740 10436
rect 3804 10372 3805 10436
rect 3739 10371 3805 10372
rect 3371 9620 3437 9621
rect 3371 9556 3372 9620
rect 3436 9556 3437 9620
rect 3371 9555 3437 9556
rect 3187 9484 3253 9485
rect 3187 9420 3188 9484
rect 3252 9420 3253 9484
rect 3187 9419 3253 9420
rect 3187 9348 3253 9349
rect 3187 9284 3188 9348
rect 3252 9284 3253 9348
rect 3187 9283 3253 9284
rect 2604 8736 2646 8954
rect 2882 8736 2924 8954
rect 2604 8672 2612 8736
rect 2676 8672 2692 8718
rect 2756 8672 2772 8718
rect 2836 8672 2852 8718
rect 2916 8672 2924 8736
rect 2604 7648 2924 8672
rect 3003 8532 3069 8533
rect 3003 8468 3004 8532
rect 3068 8468 3069 8532
rect 3003 8467 3069 8468
rect 2604 7584 2612 7648
rect 2676 7584 2692 7648
rect 2756 7584 2772 7648
rect 2836 7584 2852 7648
rect 2916 7584 2924 7648
rect 2604 6560 2924 7584
rect 2604 6496 2612 6560
rect 2676 6496 2692 6560
rect 2756 6496 2772 6560
rect 2836 6496 2852 6560
rect 2916 6496 2924 6560
rect 2604 5472 2924 6496
rect 2604 5408 2612 5472
rect 2676 5408 2692 5472
rect 2756 5408 2772 5472
rect 2836 5408 2852 5472
rect 2916 5408 2924 5472
rect 2604 4384 2924 5408
rect 3006 5269 3066 8467
rect 3003 5268 3069 5269
rect 3003 5204 3004 5268
rect 3068 5204 3069 5268
rect 3003 5203 3069 5204
rect 2604 4320 2612 4384
rect 2676 4320 2692 4384
rect 2756 4320 2772 4384
rect 2836 4320 2852 4384
rect 2916 4320 2924 4384
rect 2604 3954 2924 4320
rect 3190 4317 3250 9283
rect 3371 8396 3437 8397
rect 3371 8332 3372 8396
rect 3436 8332 3437 8396
rect 3371 8331 3437 8332
rect 3374 6901 3434 8331
rect 3558 7989 3618 10371
rect 3742 8125 3802 10371
rect 3739 8124 3805 8125
rect 3739 8060 3740 8124
rect 3804 8060 3805 8124
rect 3739 8059 3805 8060
rect 3555 7988 3621 7989
rect 3555 7924 3556 7988
rect 3620 7924 3621 7988
rect 3555 7923 3621 7924
rect 3926 7850 3986 14179
rect 4110 10845 4170 15267
rect 4294 10845 4354 15947
rect 4843 13428 4909 13429
rect 4843 13364 4844 13428
rect 4908 13364 4909 13428
rect 4843 13363 4909 13364
rect 4659 13020 4725 13021
rect 4659 12956 4660 13020
rect 4724 12956 4725 13020
rect 4659 12955 4725 12956
rect 4475 11388 4541 11389
rect 4475 11324 4476 11388
rect 4540 11324 4541 11388
rect 4475 11323 4541 11324
rect 4107 10844 4173 10845
rect 4107 10780 4108 10844
rect 4172 10780 4173 10844
rect 4107 10779 4173 10780
rect 4291 10844 4357 10845
rect 4291 10780 4292 10844
rect 4356 10780 4357 10844
rect 4291 10779 4357 10780
rect 4294 10162 4354 10422
rect 4110 10102 4354 10162
rect 4110 9077 4170 10102
rect 4291 10028 4357 10029
rect 4291 9964 4292 10028
rect 4356 9964 4357 10028
rect 4291 9963 4357 9964
rect 4107 9076 4173 9077
rect 4107 9012 4108 9076
rect 4172 9012 4173 9076
rect 4107 9011 4173 9012
rect 4107 8260 4173 8261
rect 4107 8196 4108 8260
rect 4172 8196 4173 8260
rect 4107 8195 4173 8196
rect 3742 7790 3986 7850
rect 3555 7308 3621 7309
rect 3555 7244 3556 7308
rect 3620 7244 3621 7308
rect 3555 7243 3621 7244
rect 3371 6900 3437 6901
rect 3371 6836 3372 6900
rect 3436 6836 3437 6900
rect 3371 6835 3437 6836
rect 3187 4316 3253 4317
rect 3187 4252 3188 4316
rect 3252 4252 3253 4316
rect 3187 4251 3253 4252
rect 2604 3718 2646 3954
rect 2882 3718 2924 3954
rect 2604 3296 2924 3718
rect 3371 3500 3437 3501
rect 3371 3436 3372 3500
rect 3436 3436 3437 3500
rect 3371 3435 3437 3436
rect 2604 3232 2612 3296
rect 2676 3232 2692 3296
rect 2756 3232 2772 3296
rect 2836 3232 2852 3296
rect 2916 3232 2924 3296
rect 2451 2956 2517 2957
rect 2451 2892 2452 2956
rect 2516 2892 2517 2956
rect 2451 2891 2517 2892
rect 1944 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2264 2752
rect 1347 2548 1413 2549
rect 1347 2484 1348 2548
rect 1412 2484 1413 2548
rect 1347 2483 1413 2484
rect 1944 2128 2264 2688
rect 2604 2208 2924 3232
rect 3374 2498 3434 3435
rect 3558 2685 3618 7243
rect 3742 3093 3802 7790
rect 3923 7036 3989 7037
rect 3923 6972 3924 7036
rect 3988 6972 3989 7036
rect 3923 6971 3989 6972
rect 3739 3092 3805 3093
rect 3739 3028 3740 3092
rect 3804 3028 3805 3092
rect 3739 3027 3805 3028
rect 3555 2684 3621 2685
rect 3555 2620 3556 2684
rect 3620 2620 3621 2684
rect 3555 2619 3621 2620
rect 2604 2144 2612 2208
rect 2676 2144 2692 2208
rect 2756 2144 2772 2208
rect 2836 2144 2852 2208
rect 2916 2144 2924 2208
rect 2604 2128 2924 2144
rect 3926 917 3986 6971
rect 4110 5949 4170 8195
rect 4294 6221 4354 9963
rect 4291 6220 4357 6221
rect 4291 6156 4292 6220
rect 4356 6156 4357 6220
rect 4291 6155 4357 6156
rect 4107 5948 4173 5949
rect 4107 5884 4108 5948
rect 4172 5884 4173 5948
rect 4107 5883 4173 5884
rect 4110 3501 4170 5883
rect 4478 3909 4538 11323
rect 4662 11253 4722 12955
rect 4659 11252 4725 11253
rect 4659 11188 4660 11252
rect 4724 11188 4725 11252
rect 4659 11187 4725 11188
rect 4662 9213 4722 11187
rect 4659 9212 4725 9213
rect 4659 9148 4660 9212
rect 4724 9148 4725 9212
rect 4659 9147 4725 9148
rect 4659 8940 4725 8941
rect 4659 8876 4660 8940
rect 4724 8876 4725 8940
rect 4659 8875 4725 8876
rect 4662 7853 4722 8875
rect 4659 7852 4725 7853
rect 4659 7788 4660 7852
rect 4724 7788 4725 7852
rect 4659 7787 4725 7788
rect 4659 6220 4725 6221
rect 4659 6156 4660 6220
rect 4724 6156 4725 6220
rect 4659 6155 4725 6156
rect 4475 3908 4541 3909
rect 4475 3844 4476 3908
rect 4540 3844 4541 3908
rect 4475 3843 4541 3844
rect 4107 3500 4173 3501
rect 4107 3436 4108 3500
rect 4172 3436 4173 3500
rect 4107 3435 4173 3436
rect 3923 916 3989 917
rect 3923 852 3924 916
rect 3988 852 3989 916
rect 3923 851 3989 852
rect 795 780 861 781
rect 795 716 796 780
rect 860 716 861 780
rect 795 715 861 716
rect 4662 645 4722 6155
rect 4846 5813 4906 13363
rect 5030 12341 5090 18531
rect 13859 18324 13925 18325
rect 13859 18260 13860 18324
rect 13924 18260 13925 18324
rect 13859 18259 13925 18260
rect 5763 18052 5829 18053
rect 5763 17988 5764 18052
rect 5828 17988 5829 18052
rect 5763 17987 5829 17988
rect 5395 16828 5461 16829
rect 5395 16764 5396 16828
rect 5460 16764 5461 16828
rect 5395 16763 5461 16764
rect 5398 15418 5458 16763
rect 5211 14108 5277 14109
rect 5211 14044 5212 14108
rect 5276 14044 5277 14108
rect 5211 14043 5277 14044
rect 5027 12340 5093 12341
rect 5027 12276 5028 12340
rect 5092 12276 5093 12340
rect 5027 12275 5093 12276
rect 5027 11796 5093 11797
rect 5027 11732 5028 11796
rect 5092 11732 5093 11796
rect 5027 11731 5093 11732
rect 5030 10842 5090 11731
rect 5030 10782 5136 10842
rect 5076 9621 5136 10782
rect 5214 9690 5274 14043
rect 5766 13565 5826 17987
rect 13491 17644 13557 17645
rect 13491 17580 13492 17644
rect 13556 17580 13557 17644
rect 13491 17579 13557 17580
rect 6944 16896 7264 17456
rect 6944 16832 6952 16896
rect 7016 16832 7032 16896
rect 7096 16832 7112 16896
rect 7176 16832 7192 16896
rect 7256 16832 7264 16896
rect 6315 16692 6381 16693
rect 6315 16628 6316 16692
rect 6380 16628 6381 16692
rect 6315 16627 6381 16628
rect 5763 13564 5829 13565
rect 5763 13500 5764 13564
rect 5828 13500 5829 13564
rect 5763 13499 5829 13500
rect 5947 13564 6013 13565
rect 5947 13500 5948 13564
rect 6012 13500 6013 13564
rect 5947 13499 6013 13500
rect 5950 12450 6010 13499
rect 5950 12390 6194 12450
rect 5763 12340 5829 12341
rect 5763 12276 5764 12340
rect 5828 12276 5829 12340
rect 5763 12275 5829 12276
rect 5766 12202 5826 12275
rect 5766 12142 6056 12202
rect 5579 11252 5645 11253
rect 5579 11188 5580 11252
rect 5644 11188 5645 11252
rect 5579 11187 5645 11188
rect 5395 10844 5461 10845
rect 5395 10780 5396 10844
rect 5460 10780 5461 10844
rect 5395 10779 5461 10780
rect 5398 9890 5458 10779
rect 5582 10029 5642 11187
rect 5766 10301 5826 11782
rect 5996 11522 6056 12142
rect 5950 11462 6056 11522
rect 5763 10300 5829 10301
rect 5763 10236 5764 10300
rect 5828 10236 5829 10300
rect 5763 10235 5829 10236
rect 5579 10028 5645 10029
rect 5579 9964 5580 10028
rect 5644 9964 5645 10028
rect 5579 9963 5645 9964
rect 5398 9830 5826 9890
rect 5214 9630 5458 9690
rect 5027 9620 5136 9621
rect 5027 9556 5028 9620
rect 5092 9558 5136 9620
rect 5092 9556 5093 9558
rect 5027 9555 5093 9556
rect 5027 9348 5093 9349
rect 5027 9284 5028 9348
rect 5092 9284 5093 9348
rect 5027 9283 5093 9284
rect 5211 9348 5277 9349
rect 5211 9284 5212 9348
rect 5276 9284 5277 9348
rect 5211 9283 5277 9284
rect 5030 7717 5090 9283
rect 5027 7716 5093 7717
rect 5027 7652 5028 7716
rect 5092 7652 5093 7716
rect 5027 7651 5093 7652
rect 5027 7444 5093 7445
rect 5027 7380 5028 7444
rect 5092 7380 5093 7444
rect 5027 7379 5093 7380
rect 4843 5812 4909 5813
rect 4843 5748 4844 5812
rect 4908 5748 4909 5812
rect 4843 5747 4909 5748
rect 5030 4589 5090 7379
rect 5214 4861 5274 9283
rect 5398 8669 5458 9630
rect 5766 9485 5826 9830
rect 5579 9484 5645 9485
rect 5579 9420 5580 9484
rect 5644 9420 5645 9484
rect 5579 9419 5645 9420
rect 5763 9484 5829 9485
rect 5763 9420 5764 9484
rect 5828 9420 5829 9484
rect 5763 9419 5829 9420
rect 5395 8668 5461 8669
rect 5395 8604 5396 8668
rect 5460 8604 5461 8668
rect 5395 8603 5461 8604
rect 5395 8396 5461 8397
rect 5395 8332 5396 8396
rect 5460 8332 5461 8396
rect 5395 8331 5461 8332
rect 5211 4860 5277 4861
rect 5211 4796 5212 4860
rect 5276 4796 5277 4860
rect 5211 4795 5277 4796
rect 5027 4588 5093 4589
rect 5027 4524 5028 4588
rect 5092 4524 5093 4588
rect 5027 4523 5093 4524
rect 5398 2277 5458 8331
rect 5582 5269 5642 9419
rect 5766 5813 5826 9419
rect 5950 8125 6010 11462
rect 5947 8124 6013 8125
rect 5947 8060 5948 8124
rect 6012 8060 6013 8124
rect 5947 8059 6013 8060
rect 5947 7580 6013 7581
rect 5947 7516 5948 7580
rect 6012 7516 6013 7580
rect 5947 7515 6013 7516
rect 5950 6354 6010 7515
rect 6134 7309 6194 12390
rect 6318 10709 6378 16627
rect 6944 15808 7264 16832
rect 6944 15744 6952 15808
rect 7016 15744 7032 15808
rect 7096 15744 7112 15808
rect 7176 15744 7192 15808
rect 7256 15744 7264 15808
rect 6944 14720 7264 15744
rect 7604 17440 7924 17456
rect 7604 17376 7612 17440
rect 7676 17376 7692 17440
rect 7756 17376 7772 17440
rect 7836 17376 7852 17440
rect 7916 17376 7924 17440
rect 7604 16352 7924 17376
rect 11944 16896 12264 17456
rect 11944 16832 11952 16896
rect 12016 16832 12032 16896
rect 12096 16832 12112 16896
rect 12176 16832 12192 16896
rect 12256 16832 12264 16896
rect 9075 16828 9141 16829
rect 9075 16764 9076 16828
rect 9140 16764 9141 16828
rect 9075 16763 9141 16764
rect 7604 16288 7612 16352
rect 7676 16288 7692 16352
rect 7756 16288 7772 16352
rect 7836 16288 7852 16352
rect 7916 16288 7924 16352
rect 7604 15264 7924 16288
rect 8707 15332 8773 15333
rect 8707 15268 8708 15332
rect 8772 15268 8773 15332
rect 8707 15267 8773 15268
rect 7604 15200 7612 15264
rect 7676 15200 7692 15264
rect 7756 15200 7772 15264
rect 7836 15200 7852 15264
rect 7916 15200 7924 15264
rect 7419 15196 7485 15197
rect 7419 15132 7420 15196
rect 7484 15132 7485 15196
rect 7419 15131 7485 15132
rect 7422 14789 7482 15131
rect 7419 14788 7485 14789
rect 7419 14724 7420 14788
rect 7484 14724 7485 14788
rect 7419 14723 7485 14724
rect 6944 14656 6952 14720
rect 7016 14656 7032 14720
rect 7096 14656 7112 14720
rect 7176 14656 7192 14720
rect 7256 14656 7264 14720
rect 6499 13836 6565 13837
rect 6499 13772 6500 13836
rect 6564 13772 6565 13836
rect 6499 13771 6565 13772
rect 6315 10708 6381 10709
rect 6315 10644 6316 10708
rect 6380 10644 6381 10708
rect 6315 10643 6381 10644
rect 6315 10572 6381 10573
rect 6315 10508 6316 10572
rect 6380 10508 6381 10572
rect 6315 10507 6381 10508
rect 6318 9757 6378 10507
rect 6315 9756 6381 9757
rect 6315 9692 6316 9756
rect 6380 9692 6381 9756
rect 6315 9691 6381 9692
rect 6315 9620 6381 9621
rect 6315 9556 6316 9620
rect 6380 9556 6381 9620
rect 6315 9555 6381 9556
rect 6318 9213 6378 9555
rect 6315 9212 6381 9213
rect 6315 9148 6316 9212
rect 6380 9148 6381 9212
rect 6315 9147 6381 9148
rect 6315 8940 6381 8941
rect 6315 8876 6316 8940
rect 6380 8876 6381 8940
rect 6315 8875 6381 8876
rect 6131 7308 6197 7309
rect 6131 7244 6132 7308
rect 6196 7244 6197 7308
rect 6131 7243 6197 7244
rect 5950 6294 6194 6354
rect 5947 5948 6013 5949
rect 5947 5884 5948 5948
rect 6012 5884 6013 5948
rect 5947 5883 6013 5884
rect 5763 5812 5829 5813
rect 5763 5748 5764 5812
rect 5828 5748 5829 5812
rect 5763 5747 5829 5748
rect 5579 5268 5645 5269
rect 5579 5204 5580 5268
rect 5644 5204 5645 5268
rect 5579 5203 5645 5204
rect 5950 3637 6010 5883
rect 6134 4453 6194 6294
rect 6318 4997 6378 8875
rect 6502 6765 6562 13771
rect 6944 13632 7264 14656
rect 7419 14652 7485 14653
rect 7419 14588 7420 14652
rect 7484 14588 7485 14652
rect 7419 14587 7485 14588
rect 6944 13568 6952 13632
rect 7016 13568 7032 13632
rect 7096 13568 7112 13632
rect 7176 13568 7192 13632
rect 7256 13568 7264 13632
rect 6683 13564 6749 13565
rect 6683 13500 6684 13564
rect 6748 13500 6749 13564
rect 6683 13499 6749 13500
rect 6686 8805 6746 13499
rect 6944 13294 7264 13568
rect 6944 13058 6986 13294
rect 7222 13058 7264 13294
rect 6944 12544 7264 13058
rect 6944 12480 6952 12544
rect 7016 12480 7032 12544
rect 7096 12480 7112 12544
rect 7176 12480 7192 12544
rect 7256 12480 7264 12544
rect 6944 11456 7264 12480
rect 6944 11392 6952 11456
rect 7016 11392 7032 11456
rect 7096 11392 7112 11456
rect 7176 11392 7192 11456
rect 7256 11392 7264 11456
rect 6944 10368 7264 11392
rect 7422 10981 7482 14587
rect 7604 14176 7924 15200
rect 8523 15060 8589 15061
rect 8523 14996 8524 15060
rect 8588 14996 8589 15060
rect 8523 14995 8589 14996
rect 8339 14652 8405 14653
rect 8339 14588 8340 14652
rect 8404 14588 8405 14652
rect 8339 14587 8405 14588
rect 7604 14112 7612 14176
rect 7676 14112 7692 14176
rect 7756 14112 7772 14176
rect 7836 14112 7852 14176
rect 7916 14112 7924 14176
rect 7604 13954 7924 14112
rect 7604 13718 7646 13954
rect 7882 13718 7924 13954
rect 7604 13088 7924 13718
rect 7604 13024 7612 13088
rect 7676 13024 7692 13088
rect 7756 13024 7772 13088
rect 7836 13024 7852 13088
rect 7916 13024 7924 13088
rect 7604 12000 7924 13024
rect 8155 12068 8221 12069
rect 8155 12004 8156 12068
rect 8220 12004 8221 12068
rect 8155 12003 8221 12004
rect 7604 11936 7612 12000
rect 7676 11936 7692 12000
rect 7756 11936 7772 12000
rect 7836 11936 7852 12000
rect 7916 11936 7924 12000
rect 7419 10980 7485 10981
rect 7419 10916 7420 10980
rect 7484 10916 7485 10980
rect 7419 10915 7485 10916
rect 7604 10912 7924 11936
rect 7604 10848 7612 10912
rect 7676 10848 7692 10912
rect 7756 10848 7772 10912
rect 7836 10848 7852 10912
rect 7916 10848 7924 10912
rect 7419 10844 7485 10845
rect 7419 10780 7420 10844
rect 7484 10780 7485 10844
rect 7419 10779 7485 10780
rect 6944 10304 6952 10368
rect 7016 10304 7032 10368
rect 7096 10304 7112 10368
rect 7176 10304 7192 10368
rect 7256 10304 7264 10368
rect 6944 9280 7264 10304
rect 6944 9216 6952 9280
rect 7016 9216 7032 9280
rect 7096 9216 7112 9280
rect 7176 9216 7192 9280
rect 7256 9216 7264 9280
rect 6683 8804 6749 8805
rect 6683 8740 6684 8804
rect 6748 8740 6749 8804
rect 6683 8739 6749 8740
rect 6944 8294 7264 9216
rect 6683 8260 6749 8261
rect 6683 8196 6684 8260
rect 6748 8196 6749 8260
rect 6683 8195 6749 8196
rect 6499 6764 6565 6765
rect 6499 6700 6500 6764
rect 6564 6700 6565 6764
rect 6499 6699 6565 6700
rect 6499 6220 6565 6221
rect 6499 6156 6500 6220
rect 6564 6156 6565 6220
rect 6499 6155 6565 6156
rect 6315 4996 6381 4997
rect 6315 4932 6316 4996
rect 6380 4932 6381 4996
rect 6315 4931 6381 4932
rect 6131 4452 6197 4453
rect 6131 4388 6132 4452
rect 6196 4388 6197 4452
rect 6131 4387 6197 4388
rect 6318 3909 6378 4931
rect 6315 3908 6381 3909
rect 6315 3844 6316 3908
rect 6380 3844 6381 3908
rect 6315 3843 6381 3844
rect 5947 3636 6013 3637
rect 5947 3572 5948 3636
rect 6012 3572 6013 3636
rect 5947 3571 6013 3572
rect 6502 3365 6562 6155
rect 6686 5269 6746 8195
rect 6944 8192 6986 8294
rect 7222 8192 7264 8294
rect 7422 8261 7482 10779
rect 7604 9824 7924 10848
rect 7604 9760 7612 9824
rect 7676 9760 7692 9824
rect 7756 9760 7772 9824
rect 7836 9760 7852 9824
rect 7916 9760 7924 9824
rect 7604 8954 7924 9760
rect 8158 9213 8218 12003
rect 8342 11389 8402 14587
rect 8526 13701 8586 14995
rect 8523 13700 8589 13701
rect 8523 13636 8524 13700
rect 8588 13636 8589 13700
rect 8523 13635 8589 13636
rect 8523 13156 8589 13157
rect 8523 13092 8524 13156
rect 8588 13092 8589 13156
rect 8523 13091 8589 13092
rect 8339 11388 8405 11389
rect 8339 11324 8340 11388
rect 8404 11324 8405 11388
rect 8339 11323 8405 11324
rect 8155 9212 8221 9213
rect 8155 9148 8156 9212
rect 8220 9148 8221 9212
rect 8155 9147 8221 9148
rect 7604 8736 7646 8954
rect 7882 8736 7924 8954
rect 7604 8672 7612 8736
rect 7676 8672 7692 8718
rect 7756 8672 7772 8718
rect 7836 8672 7852 8718
rect 7916 8672 7924 8736
rect 7419 8260 7485 8261
rect 7419 8196 7420 8260
rect 7484 8196 7485 8260
rect 7419 8195 7485 8196
rect 6944 8128 6952 8192
rect 7256 8128 7264 8192
rect 6944 8058 6986 8128
rect 7222 8058 7264 8128
rect 6944 7104 7264 8058
rect 6944 7040 6952 7104
rect 7016 7040 7032 7104
rect 7096 7040 7112 7104
rect 7176 7040 7192 7104
rect 7256 7040 7264 7104
rect 6944 6016 7264 7040
rect 6944 5952 6952 6016
rect 7016 5952 7032 6016
rect 7096 5952 7112 6016
rect 7176 5952 7192 6016
rect 7256 5952 7264 6016
rect 6683 5268 6749 5269
rect 6683 5204 6684 5268
rect 6748 5204 6749 5268
rect 6683 5203 6749 5204
rect 6944 4928 7264 5952
rect 7422 4997 7482 8195
rect 7604 7648 7924 8672
rect 8342 8261 8402 11323
rect 8339 8260 8405 8261
rect 8339 8196 8340 8260
rect 8404 8196 8405 8260
rect 8339 8195 8405 8196
rect 8155 7988 8221 7989
rect 8155 7924 8156 7988
rect 8220 7924 8221 7988
rect 8155 7923 8221 7924
rect 7604 7584 7612 7648
rect 7676 7584 7692 7648
rect 7756 7584 7772 7648
rect 7836 7584 7852 7648
rect 7916 7584 7924 7648
rect 7604 6560 7924 7584
rect 7604 6496 7612 6560
rect 7676 6496 7692 6560
rect 7756 6496 7772 6560
rect 7836 6496 7852 6560
rect 7916 6496 7924 6560
rect 7604 5472 7924 6496
rect 8158 6357 8218 7923
rect 8342 7853 8402 8195
rect 8339 7852 8405 7853
rect 8339 7788 8340 7852
rect 8404 7788 8405 7852
rect 8339 7787 8405 7788
rect 8339 7444 8405 7445
rect 8339 7380 8340 7444
rect 8404 7380 8405 7444
rect 8339 7379 8405 7380
rect 8155 6356 8221 6357
rect 8155 6292 8156 6356
rect 8220 6292 8221 6356
rect 8155 6291 8221 6292
rect 8155 5948 8221 5949
rect 8155 5884 8156 5948
rect 8220 5884 8221 5948
rect 8155 5883 8221 5884
rect 7604 5408 7612 5472
rect 7676 5408 7692 5472
rect 7756 5408 7772 5472
rect 7836 5408 7852 5472
rect 7916 5408 7924 5472
rect 7419 4996 7485 4997
rect 7419 4932 7420 4996
rect 7484 4932 7485 4996
rect 7419 4931 7485 4932
rect 6944 4864 6952 4928
rect 7016 4864 7032 4928
rect 7096 4864 7112 4928
rect 7176 4864 7192 4928
rect 7256 4864 7264 4928
rect 6944 3840 7264 4864
rect 7422 4453 7482 4931
rect 7419 4452 7485 4453
rect 7419 4388 7420 4452
rect 7484 4388 7485 4452
rect 7419 4387 7485 4388
rect 6944 3776 6952 3840
rect 7016 3776 7032 3840
rect 7096 3776 7112 3840
rect 7176 3776 7192 3840
rect 7256 3776 7264 3840
rect 6499 3364 6565 3365
rect 6499 3300 6500 3364
rect 6564 3300 6565 3364
rect 6499 3299 6565 3300
rect 6944 3294 7264 3776
rect 6944 3058 6986 3294
rect 7222 3058 7264 3294
rect 6944 2752 7264 3058
rect 6944 2688 6952 2752
rect 7016 2688 7032 2752
rect 7096 2688 7112 2752
rect 7176 2688 7192 2752
rect 7256 2688 7264 2752
rect 5395 2276 5461 2277
rect 5395 2212 5396 2276
rect 5460 2212 5461 2276
rect 5395 2211 5461 2212
rect 6944 2128 7264 2688
rect 7604 4384 7924 5408
rect 7604 4320 7612 4384
rect 7676 4320 7692 4384
rect 7756 4320 7772 4384
rect 7836 4320 7852 4384
rect 7916 4320 7924 4384
rect 7604 3954 7924 4320
rect 7604 3718 7646 3954
rect 7882 3718 7924 3954
rect 7604 3296 7924 3718
rect 7604 3232 7612 3296
rect 7676 3232 7692 3296
rect 7756 3232 7772 3296
rect 7836 3232 7852 3296
rect 7916 3232 7924 3296
rect 7604 2208 7924 3232
rect 8158 2685 8218 5883
rect 8342 4181 8402 7379
rect 8339 4180 8405 4181
rect 8339 4116 8340 4180
rect 8404 4116 8405 4180
rect 8339 4115 8405 4116
rect 8526 3909 8586 13091
rect 8523 3908 8589 3909
rect 8523 3844 8524 3908
rect 8588 3844 8589 3908
rect 8523 3843 8589 3844
rect 8710 2685 8770 15267
rect 9078 13157 9138 16763
rect 9443 16284 9509 16285
rect 9443 16220 9444 16284
rect 9508 16220 9509 16284
rect 9443 16219 9509 16220
rect 10731 16284 10797 16285
rect 10731 16220 10732 16284
rect 10796 16220 10797 16284
rect 10731 16219 10797 16220
rect 9259 15468 9325 15469
rect 9259 15404 9260 15468
rect 9324 15404 9325 15468
rect 9259 15403 9325 15404
rect 9075 13156 9141 13157
rect 9075 13092 9076 13156
rect 9140 13092 9141 13156
rect 9075 13091 9141 13092
rect 9075 13020 9141 13021
rect 9075 12956 9076 13020
rect 9140 12956 9141 13020
rect 9075 12955 9141 12956
rect 8891 12748 8957 12749
rect 8891 12684 8892 12748
rect 8956 12684 8957 12748
rect 8891 12683 8957 12684
rect 8894 9077 8954 12683
rect 9078 9485 9138 12955
rect 9262 12069 9322 15403
rect 9259 12068 9325 12069
rect 9259 12004 9260 12068
rect 9324 12004 9325 12068
rect 9259 12003 9325 12004
rect 9259 11388 9325 11389
rect 9259 11324 9260 11388
rect 9324 11324 9325 11388
rect 9259 11323 9325 11324
rect 9075 9484 9141 9485
rect 9075 9420 9076 9484
rect 9140 9420 9141 9484
rect 9075 9419 9141 9420
rect 8891 9076 8957 9077
rect 8891 9012 8892 9076
rect 8956 9012 8957 9076
rect 8891 9011 8957 9012
rect 8891 8804 8957 8805
rect 8891 8740 8892 8804
rect 8956 8740 8957 8804
rect 8891 8739 8957 8740
rect 8894 2685 8954 8739
rect 9078 5269 9138 9419
rect 9075 5268 9141 5269
rect 9075 5204 9076 5268
rect 9140 5204 9141 5268
rect 9075 5203 9141 5204
rect 9262 3773 9322 11323
rect 9446 10573 9506 16219
rect 10179 15876 10245 15877
rect 10179 15812 10180 15876
rect 10244 15812 10245 15876
rect 10179 15811 10245 15812
rect 9627 15196 9693 15197
rect 9627 15132 9628 15196
rect 9692 15132 9693 15196
rect 9627 15131 9693 15132
rect 9630 11389 9690 15131
rect 9811 15060 9877 15061
rect 9811 14996 9812 15060
rect 9876 14996 9877 15060
rect 9811 14995 9877 14996
rect 9814 13157 9874 14995
rect 9995 13428 10061 13429
rect 9995 13364 9996 13428
rect 10060 13364 10061 13428
rect 9995 13363 10061 13364
rect 9811 13156 9877 13157
rect 9811 13092 9812 13156
rect 9876 13092 9877 13156
rect 9811 13091 9877 13092
rect 9811 12748 9877 12749
rect 9811 12684 9812 12748
rect 9876 12684 9877 12748
rect 9811 12683 9877 12684
rect 9627 11388 9693 11389
rect 9627 11324 9628 11388
rect 9692 11324 9693 11388
rect 9627 11323 9693 11324
rect 9443 10572 9509 10573
rect 9443 10508 9444 10572
rect 9508 10508 9509 10572
rect 9443 10507 9509 10508
rect 9443 10300 9509 10301
rect 9443 10236 9444 10300
rect 9508 10236 9509 10300
rect 9443 10235 9509 10236
rect 9627 10300 9693 10301
rect 9627 10236 9628 10300
rect 9692 10236 9693 10300
rect 9627 10235 9693 10236
rect 9446 8125 9506 10235
rect 9443 8124 9509 8125
rect 9443 8060 9444 8124
rect 9508 8060 9509 8124
rect 9443 8059 9509 8060
rect 9446 7037 9506 8059
rect 9443 7036 9509 7037
rect 9443 6972 9444 7036
rect 9508 6972 9509 7036
rect 9443 6971 9509 6972
rect 9630 5133 9690 10235
rect 9814 5949 9874 12683
rect 9998 9757 10058 13363
rect 10182 11797 10242 15811
rect 10547 13428 10613 13429
rect 10547 13364 10548 13428
rect 10612 13364 10613 13428
rect 10547 13363 10613 13364
rect 10363 13292 10429 13293
rect 10363 13228 10364 13292
rect 10428 13228 10429 13292
rect 10363 13227 10429 13228
rect 10179 11796 10245 11797
rect 10179 11732 10180 11796
rect 10244 11732 10245 11796
rect 10179 11731 10245 11732
rect 10366 10301 10426 13227
rect 10550 13021 10610 13363
rect 10547 13020 10613 13021
rect 10547 12956 10548 13020
rect 10612 12956 10613 13020
rect 10547 12955 10613 12956
rect 10363 10300 10429 10301
rect 10363 10236 10364 10300
rect 10428 10236 10429 10300
rect 10363 10235 10429 10236
rect 9995 9756 10061 9757
rect 9995 9692 9996 9756
rect 10060 9754 10061 9756
rect 10060 9694 10426 9754
rect 10060 9692 10061 9694
rect 9995 9691 10061 9692
rect 10179 9212 10245 9213
rect 10179 9148 10180 9212
rect 10244 9148 10245 9212
rect 10179 9147 10245 9148
rect 9995 8532 10061 8533
rect 9995 8468 9996 8532
rect 10060 8468 10061 8532
rect 9995 8467 10061 8468
rect 9811 5948 9877 5949
rect 9811 5884 9812 5948
rect 9876 5884 9877 5948
rect 9811 5883 9877 5884
rect 9998 5541 10058 8467
rect 10182 6493 10242 9147
rect 10366 7173 10426 9694
rect 10363 7172 10429 7173
rect 10363 7108 10364 7172
rect 10428 7108 10429 7172
rect 10363 7107 10429 7108
rect 10179 6492 10245 6493
rect 10179 6428 10180 6492
rect 10244 6428 10245 6492
rect 10179 6427 10245 6428
rect 10363 6356 10429 6357
rect 10363 6292 10364 6356
rect 10428 6292 10429 6356
rect 10363 6291 10429 6292
rect 9995 5540 10061 5541
rect 9995 5476 9996 5540
rect 10060 5476 10061 5540
rect 9995 5475 10061 5476
rect 9627 5132 9693 5133
rect 9627 5068 9628 5132
rect 9692 5068 9693 5132
rect 9627 5067 9693 5068
rect 9259 3772 9325 3773
rect 9259 3708 9260 3772
rect 9324 3708 9325 3772
rect 9259 3707 9325 3708
rect 9262 3365 9322 3707
rect 9259 3364 9325 3365
rect 9259 3300 9260 3364
rect 9324 3300 9325 3364
rect 9259 3299 9325 3300
rect 8155 2684 8221 2685
rect 8155 2620 8156 2684
rect 8220 2620 8221 2684
rect 8155 2619 8221 2620
rect 8707 2684 8773 2685
rect 8707 2620 8708 2684
rect 8772 2620 8773 2684
rect 8707 2619 8773 2620
rect 8891 2684 8957 2685
rect 8891 2620 8892 2684
rect 8956 2620 8957 2684
rect 8891 2619 8957 2620
rect 10366 2549 10426 6291
rect 10363 2548 10429 2549
rect 10363 2484 10364 2548
rect 10428 2484 10429 2548
rect 10363 2483 10429 2484
rect 7604 2144 7612 2208
rect 7676 2144 7692 2208
rect 7756 2144 7772 2208
rect 7836 2144 7852 2208
rect 7916 2144 7924 2208
rect 7604 2128 7924 2144
rect 10550 1869 10610 12955
rect 10734 11253 10794 16219
rect 11944 15808 12264 16832
rect 11944 15744 11952 15808
rect 12016 15744 12032 15808
rect 12096 15744 12112 15808
rect 12176 15744 12192 15808
rect 12256 15744 12264 15808
rect 10915 15468 10981 15469
rect 10915 15404 10916 15468
rect 10980 15404 10981 15468
rect 10915 15403 10981 15404
rect 10918 12613 10978 15403
rect 11099 13292 11165 13293
rect 11099 13228 11100 13292
rect 11164 13228 11165 13292
rect 11099 13227 11165 13228
rect 10915 12612 10981 12613
rect 10915 12548 10916 12612
rect 10980 12548 10981 12612
rect 10915 12547 10981 12548
rect 10915 11796 10981 11797
rect 10915 11732 10916 11796
rect 10980 11732 10981 11796
rect 10915 11731 10981 11732
rect 10731 11252 10797 11253
rect 10731 11188 10732 11252
rect 10796 11188 10797 11252
rect 10731 11187 10797 11188
rect 10731 10844 10797 10845
rect 10731 10780 10732 10844
rect 10796 10780 10797 10844
rect 10731 10779 10797 10780
rect 10734 9077 10794 10779
rect 10731 9076 10797 9077
rect 10731 9012 10732 9076
rect 10796 9012 10797 9076
rect 10731 9011 10797 9012
rect 10731 8260 10797 8261
rect 10731 8196 10732 8260
rect 10796 8196 10797 8260
rect 10731 8195 10797 8196
rect 10734 7309 10794 8195
rect 10731 7308 10797 7309
rect 10731 7244 10732 7308
rect 10796 7244 10797 7308
rect 10731 7243 10797 7244
rect 10731 5812 10797 5813
rect 10731 5748 10732 5812
rect 10796 5748 10797 5812
rect 10731 5747 10797 5748
rect 10734 4045 10794 5747
rect 10731 4044 10797 4045
rect 10731 3980 10732 4044
rect 10796 3980 10797 4044
rect 10731 3979 10797 3980
rect 10918 2549 10978 11731
rect 11102 10709 11162 13227
rect 11286 12205 11346 15182
rect 11944 14720 12264 15744
rect 11944 14656 11952 14720
rect 12016 14656 12032 14720
rect 12096 14656 12112 14720
rect 12176 14656 12192 14720
rect 12256 14656 12264 14720
rect 11651 14516 11717 14517
rect 11651 14452 11652 14516
rect 11716 14452 11717 14516
rect 11651 14451 11717 14452
rect 11467 13700 11533 13701
rect 11467 13636 11468 13700
rect 11532 13636 11533 13700
rect 11467 13635 11533 13636
rect 11283 12204 11349 12205
rect 11283 12140 11284 12204
rect 11348 12140 11349 12204
rect 11283 12139 11349 12140
rect 11283 10844 11349 10845
rect 11283 10780 11284 10844
rect 11348 10780 11349 10844
rect 11283 10779 11349 10780
rect 11099 10708 11165 10709
rect 11099 10644 11100 10708
rect 11164 10644 11165 10708
rect 11099 10643 11165 10644
rect 11286 10570 11346 10779
rect 11102 10510 11346 10570
rect 11102 7717 11162 10510
rect 11283 9076 11349 9077
rect 11283 9012 11284 9076
rect 11348 9012 11349 9076
rect 11283 9011 11349 9012
rect 11099 7716 11165 7717
rect 11099 7652 11100 7716
rect 11164 7652 11165 7716
rect 11099 7651 11165 7652
rect 11099 7036 11165 7037
rect 11099 6972 11100 7036
rect 11164 6972 11165 7036
rect 11099 6971 11165 6972
rect 11102 4317 11162 6971
rect 11286 5541 11346 9011
rect 11470 7717 11530 13635
rect 11467 7716 11533 7717
rect 11467 7652 11468 7716
rect 11532 7652 11533 7716
rect 11467 7651 11533 7652
rect 11470 6085 11530 7651
rect 11467 6084 11533 6085
rect 11467 6020 11468 6084
rect 11532 6020 11533 6084
rect 11467 6019 11533 6020
rect 11283 5540 11349 5541
rect 11283 5476 11284 5540
rect 11348 5476 11349 5540
rect 11283 5475 11349 5476
rect 11283 5404 11349 5405
rect 11283 5340 11284 5404
rect 11348 5340 11349 5404
rect 11283 5339 11349 5340
rect 11099 4316 11165 4317
rect 11099 4252 11100 4316
rect 11164 4252 11165 4316
rect 11099 4251 11165 4252
rect 11286 3229 11346 5339
rect 11654 4045 11714 14451
rect 11944 13632 12264 14656
rect 11944 13568 11952 13632
rect 12016 13568 12032 13632
rect 12096 13568 12112 13632
rect 12176 13568 12192 13632
rect 12256 13568 12264 13632
rect 11944 13294 12264 13568
rect 11944 13058 11986 13294
rect 12222 13058 12264 13294
rect 11944 12544 12264 13058
rect 11944 12480 11952 12544
rect 12016 12480 12032 12544
rect 12096 12480 12112 12544
rect 12176 12480 12192 12544
rect 12256 12480 12264 12544
rect 11944 11456 12264 12480
rect 12604 17440 12924 17456
rect 12604 17376 12612 17440
rect 12676 17376 12692 17440
rect 12756 17376 12772 17440
rect 12836 17376 12852 17440
rect 12916 17376 12924 17440
rect 12604 16352 12924 17376
rect 13307 16828 13373 16829
rect 13307 16764 13308 16828
rect 13372 16764 13373 16828
rect 13307 16763 13373 16764
rect 12604 16288 12612 16352
rect 12676 16288 12692 16352
rect 12756 16288 12772 16352
rect 12836 16288 12852 16352
rect 12916 16288 12924 16352
rect 12604 15264 12924 16288
rect 12604 15200 12612 15264
rect 12676 15200 12692 15264
rect 12756 15200 12772 15264
rect 12836 15200 12852 15264
rect 12916 15200 12924 15264
rect 12604 14176 12924 15200
rect 13123 14788 13189 14789
rect 13123 14724 13124 14788
rect 13188 14724 13189 14788
rect 13123 14723 13189 14724
rect 12604 14112 12612 14176
rect 12676 14112 12692 14176
rect 12756 14112 12772 14176
rect 12836 14112 12852 14176
rect 12916 14112 12924 14176
rect 12604 13954 12924 14112
rect 12604 13718 12646 13954
rect 12882 13718 12924 13954
rect 12604 13088 12924 13718
rect 12604 13024 12612 13088
rect 12676 13024 12692 13088
rect 12756 13024 12772 13088
rect 12836 13024 12852 13088
rect 12916 13024 12924 13088
rect 12387 12204 12453 12205
rect 12387 12140 12388 12204
rect 12452 12140 12453 12204
rect 12387 12139 12453 12140
rect 11944 11392 11952 11456
rect 12016 11392 12032 11456
rect 12096 11392 12112 11456
rect 12176 11392 12192 11456
rect 12256 11392 12264 11456
rect 11944 10368 12264 11392
rect 11944 10304 11952 10368
rect 12016 10304 12032 10368
rect 12096 10304 12112 10368
rect 12176 10304 12192 10368
rect 12256 10304 12264 10368
rect 11944 9280 12264 10304
rect 12390 9757 12450 12139
rect 12604 12000 12924 13024
rect 12604 11936 12612 12000
rect 12676 11936 12692 12000
rect 12756 11936 12772 12000
rect 12836 11936 12852 12000
rect 12916 11936 12924 12000
rect 12604 10912 12924 11936
rect 12604 10848 12612 10912
rect 12676 10848 12692 10912
rect 12756 10848 12772 10912
rect 12836 10848 12852 10912
rect 12916 10848 12924 10912
rect 12604 9824 12924 10848
rect 12604 9760 12612 9824
rect 12676 9760 12692 9824
rect 12756 9760 12772 9824
rect 12836 9760 12852 9824
rect 12916 9760 12924 9824
rect 12387 9756 12453 9757
rect 12387 9692 12388 9756
rect 12452 9692 12453 9756
rect 12387 9691 12453 9692
rect 11944 9216 11952 9280
rect 12016 9216 12032 9280
rect 12096 9216 12112 9280
rect 12176 9216 12192 9280
rect 12256 9216 12264 9280
rect 11944 8294 12264 9216
rect 11944 8192 11986 8294
rect 12222 8192 12264 8294
rect 11944 8128 11952 8192
rect 12256 8128 12264 8192
rect 11944 8058 11986 8128
rect 12222 8058 12264 8128
rect 11944 7104 12264 8058
rect 12604 8954 12924 9760
rect 12604 8736 12646 8954
rect 12882 8736 12924 8954
rect 12604 8672 12612 8736
rect 12676 8672 12692 8718
rect 12756 8672 12772 8718
rect 12836 8672 12852 8718
rect 12916 8672 12924 8736
rect 12604 7648 12924 8672
rect 12604 7584 12612 7648
rect 12676 7584 12692 7648
rect 12756 7584 12772 7648
rect 12836 7584 12852 7648
rect 12916 7584 12924 7648
rect 12387 7172 12453 7173
rect 12387 7108 12388 7172
rect 12452 7108 12453 7172
rect 12387 7107 12453 7108
rect 11944 7040 11952 7104
rect 12016 7040 12032 7104
rect 12096 7040 12112 7104
rect 12176 7040 12192 7104
rect 12256 7040 12264 7104
rect 11944 6016 12264 7040
rect 11944 5952 11952 6016
rect 12016 5952 12032 6016
rect 12096 5952 12112 6016
rect 12176 5952 12192 6016
rect 12256 5952 12264 6016
rect 11944 4928 12264 5952
rect 12390 5405 12450 7107
rect 12604 6560 12924 7584
rect 13126 6901 13186 14723
rect 13310 12205 13370 16763
rect 13307 12204 13373 12205
rect 13307 12140 13308 12204
rect 13372 12140 13373 12204
rect 13307 12139 13373 12140
rect 13310 9893 13370 12139
rect 13494 10301 13554 17579
rect 13675 12204 13741 12205
rect 13675 12140 13676 12204
rect 13740 12140 13741 12204
rect 13675 12139 13741 12140
rect 13491 10300 13557 10301
rect 13491 10236 13492 10300
rect 13556 10236 13557 10300
rect 13491 10235 13557 10236
rect 13307 9892 13373 9893
rect 13307 9828 13308 9892
rect 13372 9828 13373 9892
rect 13307 9827 13373 9828
rect 13491 9756 13557 9757
rect 13491 9692 13492 9756
rect 13556 9692 13557 9756
rect 13491 9691 13557 9692
rect 13307 8396 13373 8397
rect 13307 8332 13308 8396
rect 13372 8332 13373 8396
rect 13307 8331 13373 8332
rect 13123 6900 13189 6901
rect 13123 6836 13124 6900
rect 13188 6836 13189 6900
rect 13123 6835 13189 6836
rect 12604 6496 12612 6560
rect 12676 6496 12692 6560
rect 12756 6496 12772 6560
rect 12836 6496 12852 6560
rect 12916 6496 12924 6560
rect 12604 5472 12924 6496
rect 12604 5408 12612 5472
rect 12676 5408 12692 5472
rect 12756 5408 12772 5472
rect 12836 5408 12852 5472
rect 12916 5408 12924 5472
rect 12387 5404 12453 5405
rect 12387 5340 12388 5404
rect 12452 5340 12453 5404
rect 12387 5339 12453 5340
rect 11944 4864 11952 4928
rect 12016 4864 12032 4928
rect 12096 4864 12112 4928
rect 12176 4864 12192 4928
rect 12256 4864 12264 4928
rect 11651 4044 11717 4045
rect 11651 3980 11652 4044
rect 11716 3980 11717 4044
rect 11651 3979 11717 3980
rect 11944 3840 12264 4864
rect 11944 3776 11952 3840
rect 12016 3776 12032 3840
rect 12096 3776 12112 3840
rect 12176 3776 12192 3840
rect 12256 3776 12264 3840
rect 11944 3294 12264 3776
rect 11283 3228 11349 3229
rect 11283 3164 11284 3228
rect 11348 3164 11349 3228
rect 11283 3163 11349 3164
rect 11944 3058 11986 3294
rect 12222 3058 12264 3294
rect 11944 2752 12264 3058
rect 11944 2688 11952 2752
rect 12016 2688 12032 2752
rect 12096 2688 12112 2752
rect 12176 2688 12192 2752
rect 12256 2688 12264 2752
rect 10915 2548 10981 2549
rect 10915 2484 10916 2548
rect 10980 2484 10981 2548
rect 10915 2483 10981 2484
rect 11944 2128 12264 2688
rect 12604 4384 12924 5408
rect 12604 4320 12612 4384
rect 12676 4320 12692 4384
rect 12756 4320 12772 4384
rect 12836 4320 12852 4384
rect 12916 4320 12924 4384
rect 12604 3954 12924 4320
rect 12604 3718 12646 3954
rect 12882 3718 12924 3954
rect 12604 3296 12924 3718
rect 12604 3232 12612 3296
rect 12676 3232 12692 3296
rect 12756 3232 12772 3296
rect 12836 3232 12852 3296
rect 12916 3232 12924 3296
rect 12604 2208 12924 3232
rect 12604 2144 12612 2208
rect 12676 2144 12692 2208
rect 12756 2144 12772 2208
rect 12836 2144 12852 2208
rect 12916 2144 12924 2208
rect 12604 2128 12924 2144
rect 10547 1868 10613 1869
rect 10547 1804 10548 1868
rect 10612 1804 10613 1868
rect 10547 1803 10613 1804
rect 4659 644 4725 645
rect 4659 580 4660 644
rect 4724 580 4725 644
rect 4659 579 4725 580
rect 13126 509 13186 6835
rect 13310 5269 13370 8331
rect 13307 5268 13373 5269
rect 13307 5204 13308 5268
rect 13372 5204 13373 5268
rect 13307 5203 13373 5204
rect 13494 4453 13554 9691
rect 13678 6493 13738 12139
rect 13862 11117 13922 18259
rect 14595 18188 14661 18189
rect 14595 18124 14596 18188
rect 14660 18124 14661 18188
rect 14595 18123 14661 18124
rect 14227 15876 14293 15877
rect 14227 15812 14228 15876
rect 14292 15812 14293 15876
rect 14227 15811 14293 15812
rect 14043 11524 14109 11525
rect 14043 11460 14044 11524
rect 14108 11460 14109 11524
rect 14043 11459 14109 11460
rect 13859 11116 13925 11117
rect 13859 11052 13860 11116
rect 13924 11052 13925 11116
rect 13859 11051 13925 11052
rect 13859 9892 13925 9893
rect 13859 9828 13860 9892
rect 13924 9828 13925 9892
rect 13859 9827 13925 9828
rect 13675 6492 13741 6493
rect 13675 6428 13676 6492
rect 13740 6428 13741 6492
rect 13675 6427 13741 6428
rect 13491 4452 13557 4453
rect 13491 4388 13492 4452
rect 13556 4388 13557 4452
rect 13491 4387 13557 4388
rect 13675 4452 13741 4453
rect 13675 4388 13676 4452
rect 13740 4388 13741 4452
rect 13675 4387 13741 4388
rect 13678 2498 13738 4387
rect 13862 3637 13922 9827
rect 14046 4045 14106 11459
rect 14230 9349 14290 15811
rect 14598 12450 14658 18123
rect 15147 17100 15213 17101
rect 15147 17036 15148 17100
rect 15212 17036 15213 17100
rect 15147 17035 15213 17036
rect 14963 14380 15029 14381
rect 14963 14316 14964 14380
rect 15028 14316 15029 14380
rect 14963 14315 15029 14316
rect 14414 12390 14658 12450
rect 14414 9349 14474 12390
rect 14779 11524 14845 11525
rect 14779 11460 14780 11524
rect 14844 11460 14845 11524
rect 14779 11459 14845 11460
rect 14595 10980 14661 10981
rect 14595 10916 14596 10980
rect 14660 10916 14661 10980
rect 14595 10915 14661 10916
rect 14227 9348 14293 9349
rect 14227 9284 14228 9348
rect 14292 9284 14293 9348
rect 14227 9283 14293 9284
rect 14411 9348 14477 9349
rect 14411 9284 14412 9348
rect 14476 9284 14477 9348
rect 14411 9283 14477 9284
rect 14043 4044 14109 4045
rect 14043 3980 14044 4044
rect 14108 3980 14109 4044
rect 14043 3979 14109 3980
rect 13859 3636 13925 3637
rect 13859 3572 13860 3636
rect 13924 3572 13925 3636
rect 13859 3571 13925 3572
rect 14414 2413 14474 9283
rect 14598 8125 14658 10915
rect 14595 8124 14661 8125
rect 14595 8060 14596 8124
rect 14660 8060 14661 8124
rect 14595 8059 14661 8060
rect 14782 4861 14842 11459
rect 14779 4860 14845 4861
rect 14779 4796 14780 4860
rect 14844 4796 14845 4860
rect 14779 4795 14845 4796
rect 14966 4181 15026 14315
rect 15150 12341 15210 17035
rect 15699 14652 15765 14653
rect 15699 14588 15700 14652
rect 15764 14588 15765 14652
rect 15699 14587 15765 14588
rect 15147 12340 15213 12341
rect 15147 12276 15148 12340
rect 15212 12276 15213 12340
rect 15147 12275 15213 12276
rect 15147 12204 15213 12205
rect 15147 12140 15148 12204
rect 15212 12140 15213 12204
rect 15147 12139 15213 12140
rect 15150 4725 15210 12139
rect 15515 10980 15581 10981
rect 15515 10916 15516 10980
rect 15580 10916 15581 10980
rect 15515 10915 15581 10916
rect 15331 10844 15397 10845
rect 15331 10780 15332 10844
rect 15396 10780 15397 10844
rect 15331 10779 15397 10780
rect 15147 4724 15213 4725
rect 15147 4660 15148 4724
rect 15212 4660 15213 4724
rect 15147 4659 15213 4660
rect 14963 4180 15029 4181
rect 14963 4116 14964 4180
rect 15028 4116 15029 4180
rect 14963 4115 15029 4116
rect 15147 4180 15213 4181
rect 15147 4116 15148 4180
rect 15212 4116 15213 4180
rect 15147 4115 15213 4116
rect 14411 2412 14477 2413
rect 14411 2348 14412 2412
rect 14476 2348 14477 2412
rect 14411 2347 14477 2348
rect 15150 1138 15210 4115
rect 15334 2005 15394 10779
rect 15518 10165 15578 10915
rect 15515 10164 15581 10165
rect 15515 10100 15516 10164
rect 15580 10100 15581 10164
rect 15515 10099 15581 10100
rect 15702 7989 15762 14587
rect 15886 11117 15946 18667
rect 16944 16896 17264 17456
rect 16944 16832 16952 16896
rect 17016 16832 17032 16896
rect 17096 16832 17112 16896
rect 17176 16832 17192 16896
rect 17256 16832 17264 16896
rect 16619 16492 16620 16542
rect 16684 16492 16685 16542
rect 16619 16491 16685 16492
rect 16944 15808 17264 16832
rect 16944 15744 16952 15808
rect 17016 15744 17032 15808
rect 17096 15744 17112 15808
rect 17176 15744 17192 15808
rect 17256 15744 17264 15808
rect 16944 14720 17264 15744
rect 16944 14656 16952 14720
rect 17016 14656 17032 14720
rect 17096 14656 17112 14720
rect 17176 14656 17192 14720
rect 17256 14656 17264 14720
rect 16619 13836 16685 13837
rect 16619 13772 16620 13836
rect 16684 13772 16685 13836
rect 16619 13771 16685 13772
rect 16251 11388 16317 11389
rect 16251 11324 16252 11388
rect 16316 11324 16317 11388
rect 16251 11323 16317 11324
rect 15883 11116 15949 11117
rect 15883 11052 15884 11116
rect 15948 11052 15949 11116
rect 15883 11051 15949 11052
rect 15883 10844 15949 10845
rect 15883 10780 15884 10844
rect 15948 10780 15949 10844
rect 15883 10779 15949 10780
rect 15886 9893 15946 10779
rect 15883 9892 15949 9893
rect 15883 9828 15884 9892
rect 15948 9828 15949 9892
rect 15883 9827 15949 9828
rect 16067 9756 16133 9757
rect 16067 9692 16068 9756
rect 16132 9692 16133 9756
rect 16067 9691 16133 9692
rect 15699 7988 15765 7989
rect 15699 7924 15700 7988
rect 15764 7924 15765 7988
rect 15699 7923 15765 7924
rect 15702 6765 15762 7923
rect 15699 6764 15765 6765
rect 15699 6700 15700 6764
rect 15764 6700 15765 6764
rect 15699 6699 15765 6700
rect 16070 4181 16130 9691
rect 16254 9621 16314 11323
rect 16435 9892 16501 9893
rect 16435 9828 16436 9892
rect 16500 9828 16501 9892
rect 16435 9827 16501 9828
rect 16251 9620 16317 9621
rect 16251 9556 16252 9620
rect 16316 9556 16317 9620
rect 16251 9555 16317 9556
rect 16251 9484 16317 9485
rect 16251 9420 16252 9484
rect 16316 9420 16317 9484
rect 16251 9419 16317 9420
rect 16067 4180 16133 4181
rect 16067 4116 16068 4180
rect 16132 4116 16133 4180
rect 16067 4115 16133 4116
rect 16254 2685 16314 9419
rect 16438 4589 16498 9827
rect 16435 4588 16501 4589
rect 16435 4524 16436 4588
rect 16500 4524 16501 4588
rect 16435 4523 16501 4524
rect 16251 2684 16317 2685
rect 16251 2620 16252 2684
rect 16316 2620 16317 2684
rect 16251 2619 16317 2620
rect 16622 2549 16682 13771
rect 16944 13632 17264 14656
rect 16944 13568 16952 13632
rect 17016 13568 17032 13632
rect 17096 13568 17112 13632
rect 17176 13568 17192 13632
rect 17256 13568 17264 13632
rect 16944 13294 17264 13568
rect 16944 13058 16986 13294
rect 17222 13058 17264 13294
rect 16944 12544 17264 13058
rect 16944 12480 16952 12544
rect 17016 12480 17032 12544
rect 17096 12480 17112 12544
rect 17176 12480 17192 12544
rect 17256 12480 17264 12544
rect 16944 11456 17264 12480
rect 16944 11392 16952 11456
rect 17016 11392 17032 11456
rect 17096 11392 17112 11456
rect 17176 11392 17192 11456
rect 17256 11392 17264 11456
rect 16944 10368 17264 11392
rect 16944 10304 16952 10368
rect 17016 10304 17032 10368
rect 17096 10304 17112 10368
rect 17176 10304 17192 10368
rect 17256 10304 17264 10368
rect 16803 9620 16869 9621
rect 16803 9556 16804 9620
rect 16868 9556 16869 9620
rect 16803 9555 16869 9556
rect 16806 3365 16866 9555
rect 16944 9280 17264 10304
rect 16944 9216 16952 9280
rect 17016 9216 17032 9280
rect 17096 9216 17112 9280
rect 17176 9216 17192 9280
rect 17256 9216 17264 9280
rect 16944 8294 17264 9216
rect 16944 8192 16986 8294
rect 17222 8192 17264 8294
rect 16944 8128 16952 8192
rect 17256 8128 17264 8192
rect 16944 8058 16986 8128
rect 17222 8058 17264 8128
rect 16944 7104 17264 8058
rect 16944 7040 16952 7104
rect 17016 7040 17032 7104
rect 17096 7040 17112 7104
rect 17176 7040 17192 7104
rect 17256 7040 17264 7104
rect 16944 6016 17264 7040
rect 16944 5952 16952 6016
rect 17016 5952 17032 6016
rect 17096 5952 17112 6016
rect 17176 5952 17192 6016
rect 17256 5952 17264 6016
rect 16944 4928 17264 5952
rect 16944 4864 16952 4928
rect 17016 4864 17032 4928
rect 17096 4864 17112 4928
rect 17176 4864 17192 4928
rect 17256 4864 17264 4928
rect 16944 3840 17264 4864
rect 16944 3776 16952 3840
rect 17016 3776 17032 3840
rect 17096 3776 17112 3840
rect 17176 3776 17192 3840
rect 17256 3776 17264 3840
rect 16803 3364 16869 3365
rect 16803 3300 16804 3364
rect 16868 3300 16869 3364
rect 16803 3299 16869 3300
rect 16944 3294 17264 3776
rect 16944 3058 16986 3294
rect 17222 3058 17264 3294
rect 16944 2752 17264 3058
rect 16944 2688 16952 2752
rect 17016 2688 17032 2752
rect 17096 2688 17112 2752
rect 17176 2688 17192 2752
rect 17256 2688 17264 2752
rect 16619 2548 16685 2549
rect 16619 2484 16620 2548
rect 16684 2484 16685 2548
rect 16619 2483 16685 2484
rect 16944 2128 17264 2688
rect 17604 17440 17924 17456
rect 17604 17376 17612 17440
rect 17676 17376 17692 17440
rect 17756 17376 17772 17440
rect 17836 17376 17852 17440
rect 17916 17376 17924 17440
rect 17604 16352 17924 17376
rect 17604 16288 17612 16352
rect 17676 16288 17692 16352
rect 17756 16288 17772 16352
rect 17836 16288 17852 16352
rect 17916 16288 17924 16352
rect 17604 15264 17924 16288
rect 18275 15468 18341 15469
rect 18275 15404 18276 15468
rect 18340 15404 18341 15468
rect 18275 15403 18341 15404
rect 17604 15200 17612 15264
rect 17676 15200 17692 15264
rect 17756 15200 17772 15264
rect 17836 15200 17852 15264
rect 17916 15200 17924 15264
rect 17604 14176 17924 15200
rect 17604 14112 17612 14176
rect 17676 14112 17692 14176
rect 17756 14112 17772 14176
rect 17836 14112 17852 14176
rect 17916 14112 17924 14176
rect 17604 13954 17924 14112
rect 17604 13718 17646 13954
rect 17882 13718 17924 13954
rect 17604 13088 17924 13718
rect 17604 13024 17612 13088
rect 17676 13024 17692 13088
rect 17756 13024 17772 13088
rect 17836 13024 17852 13088
rect 17916 13024 17924 13088
rect 17604 12000 17924 13024
rect 17604 11936 17612 12000
rect 17676 11936 17692 12000
rect 17756 11936 17772 12000
rect 17836 11936 17852 12000
rect 17916 11936 17924 12000
rect 17604 10912 17924 11936
rect 17604 10848 17612 10912
rect 17676 10848 17692 10912
rect 17756 10848 17772 10912
rect 17836 10848 17852 10912
rect 17916 10848 17924 10912
rect 17604 9824 17924 10848
rect 17604 9760 17612 9824
rect 17676 9760 17692 9824
rect 17756 9760 17772 9824
rect 17836 9760 17852 9824
rect 17916 9760 17924 9824
rect 17604 8954 17924 9760
rect 18091 9756 18157 9757
rect 18091 9692 18092 9756
rect 18156 9692 18157 9756
rect 18091 9691 18157 9692
rect 17604 8736 17646 8954
rect 17882 8736 17924 8954
rect 17604 8672 17612 8736
rect 17676 8672 17692 8718
rect 17756 8672 17772 8718
rect 17836 8672 17852 8718
rect 17916 8672 17924 8736
rect 17604 7648 17924 8672
rect 17604 7584 17612 7648
rect 17676 7584 17692 7648
rect 17756 7584 17772 7648
rect 17836 7584 17852 7648
rect 17916 7584 17924 7648
rect 17604 6560 17924 7584
rect 17604 6496 17612 6560
rect 17676 6496 17692 6560
rect 17756 6496 17772 6560
rect 17836 6496 17852 6560
rect 17916 6496 17924 6560
rect 17604 5472 17924 6496
rect 18094 5813 18154 9691
rect 18091 5812 18157 5813
rect 18091 5748 18092 5812
rect 18156 5748 18157 5812
rect 18091 5747 18157 5748
rect 18278 5677 18338 15403
rect 18827 13972 18893 13973
rect 18827 13908 18828 13972
rect 18892 13908 18893 13972
rect 18827 13907 18893 13908
rect 18643 13564 18709 13565
rect 18643 13500 18644 13564
rect 18708 13500 18709 13564
rect 18643 13499 18709 13500
rect 18459 12204 18525 12205
rect 18459 12140 18460 12204
rect 18524 12140 18525 12204
rect 18459 12139 18525 12140
rect 18275 5676 18341 5677
rect 18275 5612 18276 5676
rect 18340 5612 18341 5676
rect 18275 5611 18341 5612
rect 18462 5541 18522 12139
rect 18459 5540 18525 5541
rect 18459 5476 18460 5540
rect 18524 5476 18525 5540
rect 18459 5475 18525 5476
rect 17604 5408 17612 5472
rect 17676 5408 17692 5472
rect 17756 5408 17772 5472
rect 17836 5408 17852 5472
rect 17916 5408 17924 5472
rect 17604 4384 17924 5408
rect 17604 4320 17612 4384
rect 17676 4320 17692 4384
rect 17756 4320 17772 4384
rect 17836 4320 17852 4384
rect 17916 4320 17924 4384
rect 17604 3954 17924 4320
rect 17604 3718 17646 3954
rect 17882 3718 17924 3954
rect 17604 3296 17924 3718
rect 17604 3232 17612 3296
rect 17676 3232 17692 3296
rect 17756 3232 17772 3296
rect 17836 3232 17852 3296
rect 17916 3232 17924 3296
rect 17604 2208 17924 3232
rect 18646 2413 18706 13499
rect 18830 4045 18890 13907
rect 19011 12884 19077 12885
rect 19011 12820 19012 12884
rect 19076 12820 19077 12884
rect 19011 12819 19077 12820
rect 18827 4044 18893 4045
rect 18827 3980 18828 4044
rect 18892 3980 18893 4044
rect 18827 3979 18893 3980
rect 18643 2412 18709 2413
rect 18643 2348 18644 2412
rect 18708 2348 18709 2412
rect 18643 2347 18709 2348
rect 17604 2144 17612 2208
rect 17676 2144 17692 2208
rect 17756 2144 17772 2208
rect 17836 2144 17852 2208
rect 17916 2144 17924 2208
rect 17604 2128 17924 2144
rect 15331 2004 15397 2005
rect 15331 1940 15332 2004
rect 15396 1940 15397 2004
rect 15331 1939 15397 1940
rect 19014 1733 19074 12819
rect 19382 10165 19442 10422
rect 19379 10164 19445 10165
rect 19379 10100 19380 10164
rect 19444 10100 19445 10164
rect 19379 10099 19445 10100
rect 17907 1732 17973 1733
rect 17907 1668 17908 1732
rect 17972 1668 17973 1732
rect 17907 1667 17973 1668
rect 19011 1732 19077 1733
rect 19011 1668 19012 1732
rect 19076 1668 19077 1732
rect 19011 1667 19077 1668
rect 17910 1461 17970 1667
rect 17907 1460 17973 1461
rect 17907 1396 17908 1460
rect 17972 1396 17973 1460
rect 17907 1395 17973 1396
rect 13123 508 13189 509
rect 13123 444 13124 508
rect 13188 444 13189 508
rect 13123 443 13189 444
<< via4 >>
rect 894 16542 1130 16778
rect 1986 13058 2222 13294
rect 2646 13718 2882 13954
rect 1986 8192 2222 8294
rect 1986 8128 2016 8192
rect 2016 8128 2032 8192
rect 2032 8128 2096 8192
rect 2096 8128 2112 8192
rect 2112 8128 2176 8192
rect 2176 8128 2192 8192
rect 2192 8128 2222 8192
rect 1986 8058 2222 8128
rect 1630 7172 1866 7258
rect 1630 7108 1716 7172
rect 1716 7108 1780 7172
rect 1780 7108 1866 7172
rect 1630 7022 1866 7108
rect 1986 3058 2222 3294
rect 2646 8736 2882 8954
rect 2646 8718 2676 8736
rect 2676 8718 2692 8736
rect 2692 8718 2756 8736
rect 2756 8718 2772 8736
rect 2772 8718 2836 8736
rect 2836 8718 2852 8736
rect 2852 8718 2882 8736
rect 4160 10422 4396 10658
rect 2646 3718 2882 3954
rect 3286 2262 3522 2498
rect 1630 1052 1866 1138
rect 1630 988 1716 1052
rect 1716 988 1780 1052
rect 1780 988 1866 1052
rect 1630 902 1866 988
rect 5310 15182 5546 15418
rect 5678 11782 5914 12018
rect 6986 13058 7222 13294
rect 7646 13718 7882 13954
rect 6986 8192 7222 8294
rect 7646 8736 7882 8954
rect 7646 8718 7676 8736
rect 7676 8718 7692 8736
rect 7692 8718 7756 8736
rect 7756 8718 7772 8736
rect 7772 8718 7836 8736
rect 7836 8718 7852 8736
rect 7852 8718 7882 8736
rect 6986 8128 7016 8192
rect 7016 8128 7032 8192
rect 7032 8128 7096 8192
rect 7096 8128 7112 8192
rect 7112 8128 7176 8192
rect 7176 8128 7192 8192
rect 7192 8128 7222 8192
rect 6986 8058 7222 8128
rect 6986 3058 7222 3294
rect 7646 3718 7882 3954
rect 11198 15182 11434 15418
rect 11986 13058 12222 13294
rect 12646 13718 12882 13954
rect 11986 8192 12222 8294
rect 11986 8128 12016 8192
rect 12016 8128 12032 8192
rect 12032 8128 12096 8192
rect 12096 8128 12112 8192
rect 12112 8128 12176 8192
rect 12176 8128 12192 8192
rect 12192 8128 12222 8192
rect 11986 8058 12222 8128
rect 12646 8736 12882 8954
rect 12646 8718 12676 8736
rect 12676 8718 12692 8736
rect 12692 8718 12756 8736
rect 12756 8718 12772 8736
rect 12772 8718 12836 8736
rect 12836 8718 12852 8736
rect 12852 8718 12882 8736
rect 11986 3058 12222 3294
rect 12646 3718 12882 3954
rect 13590 2262 13826 2498
rect 16534 16556 16770 16778
rect 16534 16542 16620 16556
rect 16620 16542 16684 16556
rect 16684 16542 16770 16556
rect 16166 11932 16402 12018
rect 16166 11868 16252 11932
rect 16252 11868 16316 11932
rect 16316 11868 16402 11932
rect 16166 11782 16402 11868
rect 15614 6492 15850 6578
rect 15614 6428 15700 6492
rect 15700 6428 15764 6492
rect 15764 6428 15850 6492
rect 15614 6342 15850 6428
rect 16986 13058 17222 13294
rect 16986 8192 17222 8294
rect 16986 8128 17016 8192
rect 17016 8128 17032 8192
rect 17032 8128 17096 8192
rect 17096 8128 17112 8192
rect 17112 8128 17176 8192
rect 17176 8128 17192 8192
rect 17192 8128 17222 8192
rect 16986 8058 17222 8128
rect 16986 3058 17222 3294
rect 17646 13718 17882 13954
rect 17646 8736 17882 8954
rect 17646 8718 17676 8736
rect 17676 8718 17692 8736
rect 17692 8718 17756 8736
rect 17756 8718 17772 8736
rect 17772 8718 17836 8736
rect 17836 8718 17852 8736
rect 17852 8718 17882 8736
rect 17646 3718 17882 3954
rect 19294 10422 19530 10658
rect 15062 902 15298 1138
<< metal5 >>
rect 852 16778 16812 16820
rect 852 16542 894 16778
rect 1130 16542 16534 16778
rect 16770 16542 16812 16778
rect 852 16500 16812 16542
rect 5268 15418 11476 15460
rect 5268 15182 5310 15418
rect 5546 15182 11198 15418
rect 11434 15182 11476 15418
rect 5268 15140 11476 15182
rect 1056 13954 18908 13996
rect 1056 13718 2646 13954
rect 2882 13718 7646 13954
rect 7882 13718 12646 13954
rect 12882 13718 17646 13954
rect 17882 13718 18908 13954
rect 1056 13676 18908 13718
rect 1056 13294 18908 13336
rect 1056 13058 1986 13294
rect 2222 13058 6986 13294
rect 7222 13058 11986 13294
rect 12222 13058 16986 13294
rect 17222 13058 18908 13294
rect 1056 13016 18908 13058
rect 5636 12018 16444 12060
rect 5636 11782 5678 12018
rect 5914 11782 16166 12018
rect 16402 11782 16444 12018
rect 5636 11740 16444 11782
rect 4118 10658 19572 10700
rect 4118 10422 4160 10658
rect 4396 10422 19294 10658
rect 19530 10422 19572 10658
rect 4118 10380 19572 10422
rect 1056 8954 18908 8996
rect 1056 8718 2646 8954
rect 2882 8718 7646 8954
rect 7882 8718 12646 8954
rect 12882 8718 17646 8954
rect 17882 8718 18908 8954
rect 1056 8676 18908 8718
rect 1056 8294 18908 8336
rect 1056 8058 1986 8294
rect 2222 8058 6986 8294
rect 7222 8058 11986 8294
rect 12222 8058 16986 8294
rect 17222 8058 18908 8294
rect 1056 8016 18908 8058
rect 1588 7258 13914 7300
rect 1588 7022 1630 7258
rect 1866 7022 13914 7258
rect 1588 6980 13914 7022
rect 13594 6620 13914 6980
rect 13594 6578 15892 6620
rect 13594 6342 15614 6578
rect 15850 6342 15892 6578
rect 13594 6300 15892 6342
rect 1056 3954 18908 3996
rect 1056 3718 2646 3954
rect 2882 3718 7646 3954
rect 7882 3718 12646 3954
rect 12882 3718 17646 3954
rect 17882 3718 18908 3954
rect 1056 3676 18908 3718
rect 1056 3294 18908 3336
rect 1056 3058 1986 3294
rect 2222 3058 6986 3294
rect 7222 3058 11986 3294
rect 12222 3058 16986 3294
rect 17222 3058 18908 3294
rect 1056 3016 18908 3058
rect 3244 2498 13868 2540
rect 3244 2262 3286 2498
rect 3522 2262 13590 2498
rect 13826 2262 13868 2498
rect 3244 2220 13868 2262
rect 1588 1138 15340 1180
rect 1588 902 1630 1138
rect 1866 902 15062 1138
rect 15298 902 15340 1138
rect 1588 860 15340 902
use sky130_fd_sc_hd__clkbuf_4  _248_
timestamp 0
transform -1 0 1932 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _249_
timestamp 0
transform -1 0 11408 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _250_
timestamp 0
transform 1 0 18032 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  _251_
timestamp 0
transform -1 0 7084 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _252_
timestamp 0
transform 1 0 12052 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _253_
timestamp 0
transform -1 0 7452 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _254_
timestamp 0
transform 1 0 3956 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _255_
timestamp 0
transform 1 0 6348 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _256_
timestamp 0
transform 1 0 15088 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _257_
timestamp 0
transform -1 0 14628 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _258_
timestamp 0
transform -1 0 14996 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  _259_
timestamp 0
transform -1 0 18124 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _260_
timestamp 0
transform 1 0 6348 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _261_
timestamp 0
transform -1 0 5336 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _262_
timestamp 0
transform -1 0 6072 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _263_
timestamp 0
transform 1 0 3680 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _264_
timestamp 0
transform -1 0 6072 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _265_
timestamp 0
transform -1 0 7452 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_12  _266_
timestamp 0
transform -1 0 11500 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_4  _267_
timestamp 0
transform -1 0 10304 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_4  _268_
timestamp 0
transform -1 0 10212 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _269_
timestamp 0
transform 1 0 3036 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _270_
timestamp 0
transform 1 0 10856 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _271_
timestamp 0
transform -1 0 17020 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _272_
timestamp 0
transform 1 0 9016 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__and3_2  _273_
timestamp 0
transform -1 0 16652 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_2  _274_
timestamp 0
transform -1 0 2300 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_4  _275_
timestamp 0
transform 1 0 17112 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__a21oi_2  _276_
timestamp 0
transform -1 0 3312 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and3_4  _277_
timestamp 0
transform -1 0 2208 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _278_
timestamp 0
transform -1 0 9844 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or3_4  _279_
timestamp 0
transform 1 0 4508 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__or2b_1  _280_
timestamp 0
transform 1 0 16744 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _281_
timestamp 0
transform -1 0 6808 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _282_
timestamp 0
transform -1 0 11684 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _283_
timestamp 0
transform 1 0 2668 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _284_
timestamp 0
transform 1 0 9200 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _285_
timestamp 0
transform 1 0 11776 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _286_
timestamp 0
transform 1 0 3404 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _287_
timestamp 0
transform -1 0 7820 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _288_
timestamp 0
transform 1 0 9200 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  _289_
timestamp 0
transform -1 0 2852 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _290_
timestamp 0
transform 1 0 9568 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _291_
timestamp 0
transform 1 0 8372 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _292_
timestamp 0
transform -1 0 9568 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _293_
timestamp 0
transform 1 0 11500 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _294_
timestamp 0
transform -1 0 14168 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _295_
timestamp 0
transform 1 0 9108 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _296_
timestamp 0
transform -1 0 8924 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _297_
timestamp 0
transform 1 0 18308 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_2  _298_
timestamp 0
transform 1 0 10488 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _299_
timestamp 0
transform -1 0 10396 0 1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _300_
timestamp 0
transform -1 0 7820 0 1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__a21o_1  _301_
timestamp 0
transform 1 0 14444 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _302_
timestamp 0
transform -1 0 11408 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _303_
timestamp 0
transform 1 0 5704 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_4  _304_
timestamp 0
transform -1 0 12604 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _305_
timestamp 0
transform 1 0 1380 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _306_
timestamp 0
transform -1 0 17940 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _307_
timestamp 0
transform 1 0 14168 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _308_
timestamp 0
transform -1 0 5428 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _309_
timestamp 0
transform -1 0 7268 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  _310_
timestamp 0
transform 1 0 2852 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__and2_1  _311_
timestamp 0
transform -1 0 9292 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _312_
timestamp 0
transform -1 0 6900 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _313_
timestamp 0
transform -1 0 5520 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_2  _314_
timestamp 0
transform -1 0 8372 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__o311a_1  _315_
timestamp 0
transform -1 0 7084 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_2  _316_
timestamp 0
transform -1 0 14720 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or3_2  _317_
timestamp 0
transform 1 0 15364 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _318_
timestamp 0
transform -1 0 11960 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _319_
timestamp 0
transform 1 0 7728 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _320_
timestamp 0
transform -1 0 5704 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _321_
timestamp 0
transform -1 0 17296 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _322_
timestamp 0
transform 1 0 11500 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and4_4  _323_
timestamp 0
transform 1 0 9476 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a22oi_4  _324_
timestamp 0
transform -1 0 2944 0 1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__or3_4  _325_
timestamp 0
transform -1 0 12972 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_2  _326_
timestamp 0
transform -1 0 18584 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _327_
timestamp 0
transform -1 0 7820 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _328_
timestamp 0
transform 1 0 1748 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _329_
timestamp 0
transform 1 0 12880 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _330_
timestamp 0
transform 1 0 1380 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _331_
timestamp 0
transform -1 0 18124 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _332_
timestamp 0
transform -1 0 16008 0 1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_2  _333_
timestamp 0
transform -1 0 13616 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _334_
timestamp 0
transform 1 0 16652 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _335_
timestamp 0
transform -1 0 12696 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _336_
timestamp 0
transform 1 0 12420 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _337_
timestamp 0
transform 1 0 3956 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _338_
timestamp 0
transform -1 0 3496 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _339_
timestamp 0
transform -1 0 4692 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__buf_8  _340_
timestamp 0
transform -1 0 9384 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__a31o_1  _341_
timestamp 0
transform -1 0 16560 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__buf_6  _342_
timestamp 0
transform 1 0 10212 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _343_
timestamp 0
transform -1 0 14352 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _344_
timestamp 0
transform 1 0 6348 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _345_
timestamp 0
transform 1 0 17020 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _346_
timestamp 0
transform -1 0 9476 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _347_
timestamp 0
transform 1 0 1932 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22oi_4  _348_
timestamp 0
transform -1 0 18216 0 -1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__or3_4  _349_
timestamp 0
transform 1 0 7452 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_2  _350_
timestamp 0
transform -1 0 4416 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o21bai_2  _351_
timestamp 0
transform -1 0 7820 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _352_
timestamp 0
transform -1 0 17940 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _353_
timestamp 0
transform 1 0 8924 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _354_
timestamp 0
transform 1 0 5612 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _355_
timestamp 0
transform 1 0 15364 0 -1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_2  _356_
timestamp 0
transform 1 0 17204 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _357_
timestamp 0
transform -1 0 2944 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _358_
timestamp 0
transform 1 0 14628 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nand3b_4  _359_
timestamp 0
transform -1 0 5244 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__and3_1  _360_
timestamp 0
transform 1 0 16376 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _361_
timestamp 0
transform -1 0 12880 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _362_
timestamp 0
transform 1 0 11040 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _363_
timestamp 0
transform 1 0 11684 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _364_
timestamp 0
transform 1 0 17480 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _365_
timestamp 0
transform -1 0 12696 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _366_
timestamp 0
transform -1 0 8556 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _367_
timestamp 0
transform 1 0 5520 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _368_
timestamp 0
transform -1 0 11960 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _369_
timestamp 0
transform 1 0 18216 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _370_
timestamp 0
transform 1 0 2668 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _371_
timestamp 0
transform -1 0 18216 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _372_
timestamp 0
transform -1 0 10120 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _373_
timestamp 0
transform -1 0 17204 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__buf_6  _374_
timestamp 0
transform 1 0 2300 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _375_
timestamp 0
transform -1 0 16376 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _376_
timestamp 0
transform 1 0 14812 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _377_
timestamp 0
transform 1 0 4416 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _378_
timestamp 0
transform -1 0 11960 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _379_
timestamp 0
transform -1 0 7912 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _380_
timestamp 0
transform 1 0 12788 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _381_
timestamp 0
transform 1 0 5244 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_4  _382_
timestamp 0
transform -1 0 5336 0 -1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__a22o_4  _383_
timestamp 0
transform -1 0 7636 0 -1 5440
box -38 -48 1326 592
use sky130_fd_sc_hd__and2_4  _384_
timestamp 0
transform 1 0 5244 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _385_
timestamp 0
transform 1 0 1380 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_2  _386_
timestamp 0
transform -1 0 8372 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o21bai_4  _387_
timestamp 0
transform 1 0 5244 0 1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__nand3_4  _388_
timestamp 0
transform -1 0 3772 0 -1 4352
box -38 -48 1326 592
use sky130_fd_sc_hd__a21o_4  _389_
timestamp 0
transform -1 0 18308 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _390_
timestamp 0
transform 1 0 16652 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _391_
timestamp 0
transform 1 0 3036 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _392_
timestamp 0
transform -1 0 8464 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _393_
timestamp 0
transform 1 0 7268 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_4  _394_
timestamp 0
transform -1 0 8832 0 1 5440
box -38 -48 2062 592
use sky130_fd_sc_hd__a21o_1  _395_
timestamp 0
transform 1 0 3772 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_4  _396_
timestamp 0
transform 1 0 17296 0 -1 13056
box -38 -48 1326 592
use sky130_fd_sc_hd__a21o_1  _397_
timestamp 0
transform 1 0 4416 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and3_4  _398_
timestamp 0
transform -1 0 3404 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_2  _399_
timestamp 0
transform 1 0 1840 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _400_
timestamp 0
transform 1 0 8924 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or3_4  _401_
timestamp 0
transform 1 0 8464 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _402_
timestamp 0
transform -1 0 12420 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _403_
timestamp 0
transform 1 0 10580 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _404_
timestamp 0
transform -1 0 17020 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _405_
timestamp 0
transform 1 0 10488 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _406_
timestamp 0
transform 1 0 6440 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _407_
timestamp 0
transform 1 0 2300 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _408_
timestamp 0
transform -1 0 7636 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _409_
timestamp 0
transform -1 0 10764 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _410_
timestamp 0
transform 1 0 12604 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_2  _411_
timestamp 0
transform 1 0 4692 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _412_
timestamp 0
transform 1 0 16376 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and3_2  _413_
timestamp 0
transform -1 0 5888 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _414_
timestamp 0
transform -1 0 13340 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _415_
timestamp 0
transform -1 0 5060 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand4_4  _416_
timestamp 0
transform 1 0 3128 0 -1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__a22o_4  _417_
timestamp 0
transform -1 0 6072 0 -1 8704
box -38 -48 1326 592
use sky130_fd_sc_hd__and2_2  _418_
timestamp 0
transform 1 0 5060 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _419_
timestamp 0
transform -1 0 12052 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_2  _420_
timestamp 0
transform 1 0 17112 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _421_
timestamp 0
transform 1 0 10304 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_2  _422_
timestamp 0
transform -1 0 10396 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _423_
timestamp 0
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _424_
timestamp 0
transform -1 0 10856 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _425_
timestamp 0
transform 1 0 1564 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _426_
timestamp 0
transform -1 0 7544 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _427_
timestamp 0
transform -1 0 3036 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _428_
timestamp 0
transform 1 0 3772 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _429_
timestamp 0
transform 1 0 7912 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_2  _430_
timestamp 0
transform 1 0 4784 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _431_
timestamp 0
transform -1 0 10580 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_2  _432_
timestamp 0
transform 1 0 14076 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_2  _433_
timestamp 0
transform 1 0 4876 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and3_4  _434_
timestamp 0
transform -1 0 10028 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_2  _435_
timestamp 0
transform 1 0 2208 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a211oi_4  _436_
timestamp 0
transform -1 0 17480 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__o211a_1  _437_
timestamp 0
transform -1 0 7268 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a2111oi_4  _438_
timestamp 0
transform 1 0 16560 0 1 10880
box -38 -48 2062 592
use sky130_fd_sc_hd__or2_1  _439_
timestamp 0
transform -1 0 7912 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _440_
timestamp 0
transform 1 0 4140 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _441_
timestamp 0
transform 1 0 12328 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _442_
timestamp 0
transform -1 0 8832 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or2_4  _443_
timestamp 0
transform 1 0 14996 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _444_
timestamp 0
transform -1 0 3128 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_2  _445_
timestamp 0
transform 1 0 7452 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _446_
timestamp 0
transform 1 0 3404 0 -1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _447_
timestamp 0
transform 1 0 9568 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _448_
timestamp 0
transform 1 0 5336 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _449_
timestamp 0
transform -1 0 12972 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _450_
timestamp 0
transform -1 0 17296 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _451_
timestamp 0
transform -1 0 15824 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _452_
timestamp 0
transform 1 0 16836 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a22oi_2  _453_
timestamp 0
transform -1 0 13156 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _454_
timestamp 0
transform -1 0 11408 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _455_
timestamp 0
transform 1 0 8096 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _456_
timestamp 0
transform -1 0 13064 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _457_
timestamp 0
transform -1 0 18216 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _458_
timestamp 0
transform 1 0 5980 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _459_
timestamp 0
transform 1 0 17388 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _460_
timestamp 0
transform 1 0 12604 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _461_
timestamp 0
transform 1 0 3496 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _462_
timestamp 0
transform 1 0 14628 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _463_
timestamp 0
transform -1 0 9568 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _464_
timestamp 0
transform 1 0 16100 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _465_
timestamp 0
transform 1 0 15364 0 1 3264
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_4  _466_
timestamp 0
transform 1 0 8924 0 -1 9792
box -38 -48 1326 592
use sky130_fd_sc_hd__nand4_4  _467_
timestamp 0
transform -1 0 12052 0 1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__a22oi_2  _468_
timestamp 0
transform 1 0 6624 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__and4_1  _469_
timestamp 0
transform -1 0 11960 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_4  _470_
timestamp 0
transform -1 0 5152 0 1 6528
box -38 -48 1326 592
use sky130_fd_sc_hd__o211ai_2  _471_
timestamp 0
transform 1 0 3772 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_4  _472_
timestamp 0
transform -1 0 8096 0 1 13056
box -38 -48 1326 592
use sky130_fd_sc_hd__nand4_2  _473_
timestamp 0
transform 1 0 12144 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__a21bo_1  _474_
timestamp 0
transform -1 0 18584 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _475_
timestamp 0
transform 1 0 13156 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _476_
timestamp 0
transform -1 0 18216 0 1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__a21o_1  _477_
timestamp 0
transform -1 0 14444 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_2  _478_
timestamp 0
transform -1 0 3588 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _479_
timestamp 0
transform 1 0 7820 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _480_
timestamp 0
transform 1 0 14168 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _481_
timestamp 0
transform 1 0 5980 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _482_
timestamp 0
transform 1 0 12144 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _483_
timestamp 0
transform 1 0 11960 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _484_
timestamp 0
transform 1 0 8280 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _485_
timestamp 0
transform 1 0 11500 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__a21o_1  _486_
timestamp 0
transform -1 0 18124 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_2  _487_
timestamp 0
transform -1 0 7084 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _488_
timestamp 0
transform -1 0 12328 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _489_
timestamp 0
transform 1 0 11592 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _490_
timestamp 0
transform 1 0 10948 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a21boi_2  _491_
timestamp 0
transform 1 0 14536 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _492_
timestamp 0
transform -1 0 2116 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _493_
timestamp 0
transform -1 0 4508 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or3_4  _494_
timestamp 0
transform 1 0 4876 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _495_
timestamp 0
transform 1 0 2208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _496_
timestamp 0
transform -1 0 11224 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _497_
timestamp 0
transform -1 0 10672 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _498_
timestamp 0
transform 1 0 2852 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _499_
timestamp 0
transform 1 0 2392 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _500_
timestamp 0
transform -1 0 7912 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _501_
timestamp 0
transform -1 0 3312 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _502_
timestamp 0
transform 1 0 9200 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_4  _503_
timestamp 0
transform 1 0 13156 0 -1 15232
box -38 -48 1694 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 0
transform 1 0 16836 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 0
transform 1 0 17204 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 0
transform 1 0 5060 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 0
transform 1 0 17296 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 0
transform -1 0 18032 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 0
transform -1 0 16008 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clone7
timestamp 0
transform 1 0 8924 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_20
timestamp 0
transform 1 0 2944 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_35
timestamp 0
transform 1 0 4324 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_47
timestamp 0
transform 1 0 5428 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_55
timestamp 0
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_57
timestamp 0
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_67
timestamp 0
transform 1 0 7268 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_75
timestamp 0
transform 1 0 8004 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_83
timestamp 0
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_85
timestamp 0
transform 1 0 8924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_93
timestamp 0
transform 1 0 9660 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_103
timestamp 0
transform 1 0 10580 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_113
timestamp 0
transform 1 0 11500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_129
timestamp 0
transform 1 0 12972 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 0
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 0
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 0
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 0
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_173
timestamp 0
transform 1 0 17020 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_177
timestamp 0
transform 1 0 17388 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_9
timestamp 0
transform 1 0 1932 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_32
timestamp 0
transform 1 0 4048 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_40
timestamp 0
transform 1 0 4784 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_48
timestamp 0
transform 1 0 5520 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_65
timestamp 0
transform 1 0 7084 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_73
timestamp 0
transform 1 0 7820 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_95
timestamp 0
transform 1 0 9844 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_118
timestamp 0
transform 1 0 11960 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_122
timestamp 0
transform 1 0 12328 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_133
timestamp 0
transform 1 0 13340 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_145
timestamp 0
transform 1 0 14444 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_157
timestamp 0
transform 1 0 15548 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_165
timestamp 0
transform 1 0 16284 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_169
timestamp 0
transform 1 0 16652 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_180
timestamp 0
transform 1 0 17664 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_188
timestamp 0
transform 1 0 18400 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_9
timestamp 0
transform 1 0 1932 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_22
timestamp 0
transform 1 0 3128 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_29
timestamp 0
transform 1 0 3772 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_39
timestamp 0
transform 1 0 4692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_51
timestamp 0
transform 1 0 5796 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_58
timestamp 0
transform 1 0 6440 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_70
timestamp 0
transform 1 0 7544 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_91
timestamp 0
transform 1 0 9476 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_103
timestamp 0
transform 1 0 10580 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_115
timestamp 0
transform 1 0 11684 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_130
timestamp 0
transform 1 0 13064 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_138
timestamp 0
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 0
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_153
timestamp 0
transform 1 0 15180 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_172
timestamp 0
transform 1 0 16928 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_186
timestamp 0
transform 1 0 18216 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_3
timestamp 0
transform 1 0 1380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_7
timestamp 0
transform 1 0 1748 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_52
timestamp 0
transform 1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 0
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_69
timestamp 0
transform 1 0 7452 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_77
timestamp 0
transform 1 0 8188 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_90
timestamp 0
transform 1 0 9384 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_98
timestamp 0
transform 1 0 10120 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_110
timestamp 0
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_113
timestamp 0
transform 1 0 11500 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_126
timestamp 0
transform 1 0 12696 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_138
timestamp 0
transform 1 0 13800 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_150
timestamp 0
transform 1 0 14904 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_162
timestamp 0
transform 1 0 16008 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_173
timestamp 0
transform 1 0 17020 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_185
timestamp 0
transform 1 0 18124 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_20
timestamp 0
transform 1 0 2944 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_36
timestamp 0
transform 1 0 4416 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_52
timestamp 0
transform 1 0 5888 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_74
timestamp 0
transform 1 0 7912 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_82
timestamp 0
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 0
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_119
timestamp 0
transform 1 0 12052 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_131
timestamp 0
transform 1 0 13156 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 0
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_141
timestamp 0
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_150
timestamp 0
transform 1 0 14904 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_158
timestamp 0
transform 1 0 15640 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_170
timestamp 0
transform 1 0 16744 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_182
timestamp 0
transform 1 0 17848 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 0
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_15
timestamp 0
transform 1 0 2484 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_21
timestamp 0
transform 1 0 3036 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_47
timestamp 0
transform 1 0 5428 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 0
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_79
timestamp 0
transform 1 0 8372 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_83
timestamp 0
transform 1 0 8740 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_89
timestamp 0
transform 1 0 9292 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_101
timestamp 0
transform 1 0 10396 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_109
timestamp 0
transform 1 0 11132 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_113
timestamp 0
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_120
timestamp 0
transform 1 0 12144 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_126
timestamp 0
transform 1 0 12696 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_138
timestamp 0
transform 1 0 13800 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_150
timestamp 0
transform 1 0 14904 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_154
timestamp 0
transform 1 0 15272 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_174
timestamp 0
transform 1 0 17112 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_180
timestamp 0
transform 1 0 17664 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_186
timestamp 0
transform 1 0 18216 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_3
timestamp 0
transform 1 0 1380 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_11
timestamp 0
transform 1 0 2116 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_18
timestamp 0
transform 1 0 2760 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_36
timestamp 0
transform 1 0 4416 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_48
timestamp 0
transform 1 0 5520 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_54
timestamp 0
transform 1 0 6072 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_92
timestamp 0
transform 1 0 9568 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_100
timestamp 0
transform 1 0 10304 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_106
timestamp 0
transform 1 0 10856 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_115
timestamp 0
transform 1 0 11684 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_125
timestamp 0
transform 1 0 12604 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_137
timestamp 0
transform 1 0 13708 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_141
timestamp 0
transform 1 0 14076 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_162
timestamp 0
transform 1 0 16008 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_173
timestamp 0
transform 1 0 17020 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_177
timestamp 0
transform 1 0 17388 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_185
timestamp 0
transform 1 0 18124 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_189
timestamp 0
transform 1 0 18492 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 0
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_15
timestamp 0
transform 1 0 2484 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_23
timestamp 0
transform 1 0 3220 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_37
timestamp 0
transform 1 0 4508 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 0
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 0
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 0
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_69
timestamp 0
transform 1 0 7452 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_80
timestamp 0
transform 1 0 8464 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_88
timestamp 0
transform 1 0 9200 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_100
timestamp 0
transform 1 0 10304 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_113
timestamp 0
transform 1 0 11500 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_119
timestamp 0
transform 1 0 12052 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_123
timestamp 0
transform 1 0 12420 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_135
timestamp 0
transform 1 0 13524 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_147
timestamp 0
transform 1 0 14628 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_159
timestamp 0
transform 1 0 15732 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 0
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 0
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_181
timestamp 0
transform 1 0 17756 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_189
timestamp 0
transform 1 0 18492 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_7
timestamp 0
transform 1 0 1748 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_19
timestamp 0
transform 1 0 2852 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 0
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_29
timestamp 0
transform 1 0 3772 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_44
timestamp 0
transform 1 0 5152 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_56
timestamp 0
transform 1 0 6256 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_80
timestamp 0
transform 1 0 8464 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 0
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 0
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 0
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_121
timestamp 0
transform 1 0 12236 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_131
timestamp 0
transform 1 0 13156 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 0
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 0
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 0
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_165
timestamp 0
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_177
timestamp 0
transform 1 0 17388 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_185
timestamp 0
transform 1 0 18124 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 0
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 0
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_27
timestamp 0
transform 1 0 3588 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_33
timestamp 0
transform 1 0 4140 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_44
timestamp 0
transform 1 0 5152 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 0
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_91
timestamp 0
transform 1 0 9476 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_101
timestamp 0
transform 1 0 10396 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_105
timestamp 0
transform 1 0 10764 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_110
timestamp 0
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_118
timestamp 0
transform 1 0 11960 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_130
timestamp 0
transform 1 0 13064 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_151
timestamp 0
transform 1 0 14996 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_163
timestamp 0
transform 1 0 16100 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 0
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_169
timestamp 0
transform 1 0 16652 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_176
timestamp 0
transform 1 0 17296 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_188
timestamp 0
transform 1 0 18400 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_9
timestamp 0
transform 1 0 1932 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_20
timestamp 0
transform 1 0 2944 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_29
timestamp 0
transform 1 0 3772 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_33
timestamp 0
transform 1 0 4140 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_38
timestamp 0
transform 1 0 4600 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_50
timestamp 0
transform 1 0 5704 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_54
timestamp 0
transform 1 0 6072 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_58
timestamp 0
transform 1 0 6440 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_67
timestamp 0
transform 1 0 7268 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_79
timestamp 0
transform 1 0 8372 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 0
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_85
timestamp 0
transform 1 0 8924 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_95
timestamp 0
transform 1 0 9844 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_107
timestamp 0
transform 1 0 10948 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_119
timestamp 0
transform 1 0 12052 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_127
timestamp 0
transform 1 0 12788 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp 0
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 0
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_141
timestamp 0
transform 1 0 14076 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_149
timestamp 0
transform 1 0 14812 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_166
timestamp 0
transform 1 0 16376 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_174
timestamp 0
transform 1 0 17112 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_185
timestamp 0
transform 1 0 18124 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_189
timestamp 0
transform 1 0 18492 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_3
timestamp 0
transform 1 0 1380 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_38
timestamp 0
transform 1 0 4600 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_54
timestamp 0
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 0
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_81
timestamp 0
transform 1 0 8556 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_87
timestamp 0
transform 1 0 9108 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_104
timestamp 0
transform 1 0 10672 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 0
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 0
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_137
timestamp 0
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_149
timestamp 0
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_161
timestamp 0
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 0
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_176
timestamp 0
transform 1 0 17296 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_188
timestamp 0
transform 1 0 18400 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_15
timestamp 0
transform 1 0 2484 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_38
timestamp 0
transform 1 0 4600 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_47
timestamp 0
transform 1 0 5428 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_59
timestamp 0
transform 1 0 6532 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_67
timestamp 0
transform 1 0 7268 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_82
timestamp 0
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_110
timestamp 0
transform 1 0 11224 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_122
timestamp 0
transform 1 0 12328 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_134
timestamp 0
transform 1 0 13432 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 0
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_153
timestamp 0
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_165
timestamp 0
transform 1 0 16284 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_175
timestamp 0
transform 1 0 17204 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_181
timestamp 0
transform 1 0 17756 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_185
timestamp 0
transform 1 0 18124 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_3
timestamp 0
transform 1 0 1380 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_11
timestamp 0
transform 1 0 2116 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_25
timestamp 0
transform 1 0 3404 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_42
timestamp 0
transform 1 0 4968 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_54
timestamp 0
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_57
timestamp 0
transform 1 0 6348 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_63
timestamp 0
transform 1 0 6900 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_73
timestamp 0
transform 1 0 7820 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_108
timestamp 0
transform 1 0 11040 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_113
timestamp 0
transform 1 0 11500 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_125
timestamp 0
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_137
timestamp 0
transform 1 0 13708 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_151
timestamp 0
transform 1 0 14996 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_163
timestamp 0
transform 1 0 16100 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_167
timestamp 0
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_173
timestamp 0
transform 1 0 17020 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_3
timestamp 0
transform 1 0 1380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 0
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_29
timestamp 0
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_36
timestamp 0
transform 1 0 4416 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_48
timestamp 0
transform 1 0 5520 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_60
timestamp 0
transform 1 0 6624 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_64
timestamp 0
transform 1 0 6992 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_74
timestamp 0
transform 1 0 7912 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_82
timestamp 0
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_85
timestamp 0
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_97
timestamp 0
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_109
timestamp 0
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_121
timestamp 0
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_133
timestamp 0
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 0
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_141
timestamp 0
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_153
timestamp 0
transform 1 0 15180 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_161
timestamp 0
transform 1 0 15916 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 0
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_15
timestamp 0
transform 1 0 2484 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_28
timestamp 0
transform 1 0 3680 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_39
timestamp 0
transform 1 0 4692 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_45
timestamp 0
transform 1 0 5244 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_54
timestamp 0
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_70
timestamp 0
transform 1 0 7544 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_82
timestamp 0
transform 1 0 8648 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_94
timestamp 0
transform 1 0 9752 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_106
timestamp 0
transform 1 0 10856 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_118
timestamp 0
transform 1 0 11960 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_130
timestamp 0
transform 1 0 13064 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_136
timestamp 0
transform 1 0 13616 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_144
timestamp 0
transform 1 0 14352 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_167
timestamp 0
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_169
timestamp 0
transform 1 0 16652 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_176
timestamp 0
transform 1 0 17296 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_9
timestamp 0
transform 1 0 1932 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_21
timestamp 0
transform 1 0 3036 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 0
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_52
timestamp 0
transform 1 0 5888 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_56
timestamp 0
transform 1 0 6256 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_64
timestamp 0
transform 1 0 6992 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_73
timestamp 0
transform 1 0 7820 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_81
timestamp 0
transform 1 0 8556 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_85
timestamp 0
transform 1 0 8924 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_101
timestamp 0
transform 1 0 10396 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_109
timestamp 0
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_121
timestamp 0
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_133
timestamp 0
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 0
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_141
timestamp 0
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_153
timestamp 0
transform 1 0 15180 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_159
timestamp 0
transform 1 0 15732 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_162
timestamp 0
transform 1 0 16008 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_3
timestamp 0
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_10
timestamp 0
transform 1 0 2024 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_18
timestamp 0
transform 1 0 2760 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_35
timestamp 0
transform 1 0 4324 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_50
timestamp 0
transform 1 0 5704 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_65
timestamp 0
transform 1 0 7084 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_81
timestamp 0
transform 1 0 8556 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_89
timestamp 0
transform 1 0 9292 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_95
timestamp 0
transform 1 0 9844 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 0
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_113
timestamp 0
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_125
timestamp 0
transform 1 0 12604 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_133
timestamp 0
transform 1 0 13340 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_149
timestamp 0
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_161
timestamp 0
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_167
timestamp 0
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_169
timestamp 0
transform 1 0 16652 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_187
timestamp 0
transform 1 0 18308 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_3
timestamp 0
transform 1 0 1380 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_11
timestamp 0
transform 1 0 2116 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_22
timestamp 0
transform 1 0 3128 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_39
timestamp 0
transform 1 0 4692 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_54
timestamp 0
transform 1 0 6072 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_66
timestamp 0
transform 1 0 7176 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_78
timestamp 0
transform 1 0 8280 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_85
timestamp 0
transform 1 0 8924 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_91
timestamp 0
transform 1 0 9476 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_106
timestamp 0
transform 1 0 10856 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_118
timestamp 0
transform 1 0 11960 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_135
timestamp 0
transform 1 0 13524 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 0
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_148
timestamp 0
transform 1 0 14720 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_160
timestamp 0
transform 1 0 15824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_3
timestamp 0
transform 1 0 1380 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_11
timestamp 0
transform 1 0 2116 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_32
timestamp 0
transform 1 0 4048 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_48
timestamp 0
transform 1 0 5520 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_57
timestamp 0
transform 1 0 6348 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_73
timestamp 0
transform 1 0 7820 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_85
timestamp 0
transform 1 0 8924 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_93
timestamp 0
transform 1 0 9660 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_109
timestamp 0
transform 1 0 11132 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_128
timestamp 0
transform 1 0 12880 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_140
timestamp 0
transform 1 0 13984 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_152
timestamp 0
transform 1 0 15088 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_160
timestamp 0
transform 1 0 15824 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_169
timestamp 0
transform 1 0 16652 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_175
timestamp 0
transform 1 0 17204 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_3
timestamp 0
transform 1 0 1380 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_11
timestamp 0
transform 1 0 2116 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_24
timestamp 0
transform 1 0 3312 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 0
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_41
timestamp 0
transform 1 0 4876 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_60
timestamp 0
transform 1 0 6624 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_76
timestamp 0
transform 1 0 8096 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_85
timestamp 0
transform 1 0 8924 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_97
timestamp 0
transform 1 0 10028 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_105
timestamp 0
transform 1 0 10764 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_115
timestamp 0
transform 1 0 11684 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_123
timestamp 0
transform 1 0 12420 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_129
timestamp 0
transform 1 0 12972 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_137
timestamp 0
transform 1 0 13708 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_141
timestamp 0
transform 1 0 14076 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_149
timestamp 0
transform 1 0 14812 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_157
timestamp 0
transform 1 0 15548 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_169
timestamp 0
transform 1 0 16652 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_9
timestamp 0
transform 1 0 1932 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_24
timestamp 0
transform 1 0 3312 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_36
timestamp 0
transform 1 0 4416 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_42
timestamp 0
transform 1 0 4968 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_74
timestamp 0
transform 1 0 7912 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_80
timestamp 0
transform 1 0 8464 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_89
timestamp 0
transform 1 0 9292 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_101
timestamp 0
transform 1 0 10396 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_109
timestamp 0
transform 1 0 11132 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_113
timestamp 0
transform 1 0 11500 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_119
timestamp 0
transform 1 0 12052 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_130
timestamp 0
transform 1 0 13064 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_142
timestamp 0
transform 1 0 14168 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_154
timestamp 0
transform 1 0 15272 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_166
timestamp 0
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_169
timestamp 0
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_181
timestamp 0
transform 1 0 17756 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_189
timestamp 0
transform 1 0 18492 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_3
timestamp 0
transform 1 0 1380 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_14
timestamp 0
transform 1 0 2392 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_26
timestamp 0
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_29
timestamp 0
transform 1 0 3772 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_37
timestamp 0
transform 1 0 4508 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_43
timestamp 0
transform 1 0 5060 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_55
timestamp 0
transform 1 0 6164 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_67
timestamp 0
transform 1 0 7268 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_79
timestamp 0
transform 1 0 8372 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 0
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_85
timestamp 0
transform 1 0 8924 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_95
timestamp 0
transform 1 0 9844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_107
timestamp 0
transform 1 0 10948 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_134
timestamp 0
transform 1 0 13432 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_149
timestamp 0
transform 1 0 14812 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_161
timestamp 0
transform 1 0 15916 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_173
timestamp 0
transform 1 0 17020 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_185
timestamp 0
transform 1 0 18124 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_189
timestamp 0
transform 1 0 18492 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_9
timestamp 0
transform 1 0 1932 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_21
timestamp 0
transform 1 0 3036 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_33
timestamp 0
transform 1 0 4140 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_46
timestamp 0
transform 1 0 5336 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_54
timestamp 0
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_57
timestamp 0
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_69
timestamp 0
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_81
timestamp 0
transform 1 0 8556 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_89
timestamp 0
transform 1 0 9292 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_99
timestamp 0
transform 1 0 10212 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_108
timestamp 0
transform 1 0 11040 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_118
timestamp 0
transform 1 0 11960 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_149
timestamp 0
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_161
timestamp 0
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_167
timestamp 0
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_186
timestamp 0
transform 1 0 18216 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 0
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp 0
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 0
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_35
timestamp 0
transform 1 0 4324 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_49
timestamp 0
transform 1 0 5612 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_55
timestamp 0
transform 1 0 6164 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_65
timestamp 0
transform 1 0 7084 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_92
timestamp 0
transform 1 0 9568 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_100
timestamp 0
transform 1 0 10304 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_119
timestamp 0
transform 1 0 12052 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_134
timestamp 0
transform 1 0 13432 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_141
timestamp 0
transform 1 0 14076 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_155
timestamp 0
transform 1 0 15364 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_167
timestamp 0
transform 1 0 16468 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_179
timestamp 0
transform 1 0 17572 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_187
timestamp 0
transform 1 0 18308 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 0
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_15
timestamp 0
transform 1 0 2484 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_24
timestamp 0
transform 1 0 3312 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_36
timestamp 0
transform 1 0 4416 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_48
timestamp 0
transform 1 0 5520 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_65
timestamp 0
transform 1 0 7084 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_77
timestamp 0
transform 1 0 8188 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_89
timestamp 0
transform 1 0 9292 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_101
timestamp 0
transform 1 0 10396 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_109
timestamp 0
transform 1 0 11132 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_113
timestamp 0
transform 1 0 11500 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_119
timestamp 0
transform 1 0 12052 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_123
timestamp 0
transform 1 0 12420 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_129
timestamp 0
transform 1 0 12972 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_141
timestamp 0
transform 1 0 14076 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_153
timestamp 0
transform 1 0 15180 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_165
timestamp 0
transform 1 0 16284 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_169
timestamp 0
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_173
timestamp 0
transform 1 0 17020 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_185
timestamp 0
transform 1 0 18124 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_189
timestamp 0
transform 1 0 18492 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_13
timestamp 0
transform 1 0 2300 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_25
timestamp 0
transform 1 0 3404 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 0
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_41
timestamp 0
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_53
timestamp 0
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_65
timestamp 0
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_77
timestamp 0
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 0
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_85
timestamp 0
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_97
timestamp 0
transform 1 0 10028 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_105
timestamp 0
transform 1 0 10764 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_112
timestamp 0
transform 1 0 11408 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_124
timestamp 0
transform 1 0 12512 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_136
timestamp 0
transform 1 0 13616 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_141
timestamp 0
transform 1 0 14076 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_145
timestamp 0
transform 1 0 14444 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_155
timestamp 0
transform 1 0 15364 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_163
timestamp 0
transform 1 0 16100 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_175
timestamp 0
transform 1 0 17204 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_181
timestamp 0
transform 1 0 17756 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_184
timestamp 0
transform 1 0 18032 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_3
timestamp 0
transform 1 0 1380 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_19
timestamp 0
transform 1 0 2852 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_27
timestamp 0
transform 1 0 3588 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_35
timestamp 0
transform 1 0 4324 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_43
timestamp 0
transform 1 0 5060 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_52
timestamp 0
transform 1 0 5888 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_63
timestamp 0
transform 1 0 6900 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_75
timestamp 0
transform 1 0 8004 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_83
timestamp 0
transform 1 0 8740 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_95
timestamp 0
transform 1 0 9844 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_107
timestamp 0
transform 1 0 10948 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_126
timestamp 0
transform 1 0 12696 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_138
timestamp 0
transform 1 0 13800 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_145
timestamp 0
transform 1 0 14444 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_157
timestamp 0
transform 1 0 15548 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_169
timestamp 0
transform 1 0 16652 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_175
timestamp 0
transform 1 0 17204 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_178
timestamp 0
transform 1 0 17480 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_4  input1
timestamp 0
transform 1 0 2300 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input2
timestamp 0
transform 1 0 1380 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input3
timestamp 0
transform 1 0 1380 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input4
timestamp 0
transform 1 0 1380 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input5
timestamp 0
transform 1 0 1932 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 0
transform 1 0 1380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input7
timestamp 0
transform 1 0 1380 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input8
timestamp 0
transform 1 0 2576 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input9
timestamp 0
transform -1 0 18584 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  input10
timestamp 0
transform -1 0 16560 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  input11
timestamp 0
transform 1 0 14076 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input12
timestamp 0
transform 1 0 11040 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 0
transform 1 0 9476 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input14
timestamp 0
transform 1 0 6348 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input15
timestamp 0
transform 1 0 3772 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 0
transform 1 0 1932 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input17
timestamp 0
transform 1 0 16652 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input18
timestamp 0
transform 1 0 10028 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input19
timestamp 0
transform 1 0 3772 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  max_cap28
timestamp 0
transform 1 0 13248 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output20
timestamp 0
transform 1 0 17664 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp 0
transform 1 0 18216 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp 0
transform 1 0 18216 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 0
transform 1 0 16192 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 0
transform 1 0 18216 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp 0
transform 1 0 18216 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 0
transform 1 0 18216 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  output27
timestamp 0
transform 1 0 17480 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_28
timestamp 0
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 0
transform -1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_29
timestamp 0
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 0
transform -1 0 18860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_30
timestamp 0
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 0
transform -1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_31
timestamp 0
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 0
transform -1 0 18860 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_32
timestamp 0
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 0
transform -1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_33
timestamp 0
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 0
transform -1 0 18860 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_34
timestamp 0
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 0
transform -1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_35
timestamp 0
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 0
transform -1 0 18860 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_36
timestamp 0
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 0
transform -1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_37
timestamp 0
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 0
transform -1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_38
timestamp 0
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 0
transform -1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_39
timestamp 0
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 0
transform -1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_40
timestamp 0
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 0
transform -1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_41
timestamp 0
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 0
transform -1 0 18860 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_42
timestamp 0
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 0
transform -1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_43
timestamp 0
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 0
transform -1 0 18860 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_44
timestamp 0
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 0
transform -1 0 18860 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_45
timestamp 0
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 0
transform -1 0 18860 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_46
timestamp 0
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 0
transform -1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_47
timestamp 0
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 0
transform -1 0 18860 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_48
timestamp 0
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 0
transform -1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_49
timestamp 0
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 0
transform -1 0 18860 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_50
timestamp 0
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 0
transform -1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_51
timestamp 0
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 0
transform -1 0 18860 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_52
timestamp 0
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 0
transform -1 0 18860 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_53
timestamp 0
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 0
transform -1 0 18860 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_54
timestamp 0
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 0
transform -1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_55
timestamp 0
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 0
transform -1 0 18860 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  rebuffer1
timestamp 0
transform -1 0 3680 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer2
timestamp 0
transform 1 0 3036 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  rebuffer3
timestamp 0
transform 1 0 4232 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  rebuffer4
timestamp 0
transform 1 0 4232 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  rebuffer5
timestamp 0
transform 1 0 16652 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  rebuffer6
timestamp 0
transform 1 0 16836 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  rebuffer8
timestamp 0
transform -1 0 4600 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer9
timestamp 0
transform 1 0 3772 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  rebuffer10
timestamp 0
transform 1 0 2484 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  rebuffer11
timestamp 0
transform 1 0 5244 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  rebuffer12
timestamp 0
transform -1 0 13432 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer13
timestamp 0
transform 1 0 2024 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_56
timestamp 0
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_57
timestamp 0
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_58
timestamp 0
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_59
timestamp 0
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_60
timestamp 0
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_61
timestamp 0
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_62
timestamp 0
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_63
timestamp 0
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_64
timestamp 0
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_65
timestamp 0
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_66
timestamp 0
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_67
timestamp 0
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_68
timestamp 0
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_69
timestamp 0
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_70
timestamp 0
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_71
timestamp 0
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_72
timestamp 0
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_73
timestamp 0
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_74
timestamp 0
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_75
timestamp 0
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_76
timestamp 0
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_77
timestamp 0
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_78
timestamp 0
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_79
timestamp 0
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_80
timestamp 0
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_81
timestamp 0
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_82
timestamp 0
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_83
timestamp 0
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_84
timestamp 0
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_85
timestamp 0
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_86
timestamp 0
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_87
timestamp 0
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_88
timestamp 0
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_89
timestamp 0
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_90
timestamp 0
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_91
timestamp 0
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_92
timestamp 0
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_93
timestamp 0
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_94
timestamp 0
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_95
timestamp 0
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_96
timestamp 0
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_97
timestamp 0
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_98
timestamp 0
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_99
timestamp 0
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_100
timestamp 0
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_101
timestamp 0
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_102
timestamp 0
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_103
timestamp 0
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_104
timestamp 0
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_105
timestamp 0
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_106
timestamp 0
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_107
timestamp 0
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_108
timestamp 0
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_109
timestamp 0
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_110
timestamp 0
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_111
timestamp 0
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_112
timestamp 0
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_113
timestamp 0
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_114
timestamp 0
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_115
timestamp 0
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_116
timestamp 0
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_117
timestamp 0
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_118
timestamp 0
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_119
timestamp 0
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_120
timestamp 0
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_121
timestamp 0
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_122
timestamp 0
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_123
timestamp 0
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_124
timestamp 0
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_125
timestamp 0
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_126
timestamp 0
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_127
timestamp 0
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_128
timestamp 0
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_129
timestamp 0
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_130
timestamp 0
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_131
timestamp 0
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_132
timestamp 0
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_133
timestamp 0
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_134
timestamp 0
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_135
timestamp 0
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_136
timestamp 0
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_137
timestamp 0
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_138
timestamp 0
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_139
timestamp 0
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_140
timestamp 0
transform 1 0 3680 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_141
timestamp 0
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_142
timestamp 0
transform 1 0 8832 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_143
timestamp 0
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_144
timestamp 0
transform 1 0 13984 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_145
timestamp 0
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
<< labels >>
rlabel metal1 s 9982 17408 9982 17408 4 VGND
rlabel metal1 s 9982 16864 9982 16864 4 VPWR
rlabel metal2 s 2990 17901 2990 17901 4 A[0]
rlabel metal3 s 1096 16116 1096 16116 4 A[1]
rlabel metal3 s 1096 13668 1096 13668 4 A[2]
rlabel metal3 s 1050 11220 1050 11220 4 A[3]
rlabel metal3 s 1326 8772 1326 8772 4 A[4]
rlabel metal3 s 1096 6324 1096 6324 4 A[5]
rlabel metal3 s 1050 3876 1050 3876 4 A[6]
rlabel metal3 s 1556 1428 1556 1428 4 A[7]
rlabel metal1 s 18584 17170 18584 17170 4 B[0]
rlabel metal1 s 16284 17170 16284 17170 4 B[1]
rlabel metal1 s 13892 17170 13892 17170 4 B[2]
rlabel metal1 s 11132 17170 11132 17170 4 B[3]
rlabel metal1 s 9154 17238 9154 17238 4 B[4]
rlabel metal1 s 6348 17238 6348 17238 4 B[5]
rlabel metal1 s 3818 17238 3818 17238 4 B[6]
rlabel metal1 s 1656 16558 1656 16558 4 B[7]
rlabel metal1 s 4554 13702 4554 13702 4 _000_
rlabel metal1 s 16882 3706 16882 3706 4 _001_
rlabel metal2 s 13018 1836 13018 1836 4 _002_
rlabel metal4 s 15548 10540 15548 10540 4 _003_
rlabel metal3 s 15019 2652 15019 2652 4 _004_
rlabel metal1 s 1564 15130 1564 15130 4 _005_
rlabel metal1 s 1518 15062 1518 15062 4 _006_
rlabel metal2 s 2254 14518 2254 14518 4 _007_
rlabel metal1 s 1610 14960 1610 14960 4 _008_
rlabel metal1 s 13340 7990 13340 7990 4 _009_
rlabel metal2 s 4002 16252 4002 16252 4 _010_
rlabel metal1 s 16054 13702 16054 13702 4 _011_
rlabel metal2 s 14858 6324 14858 6324 4 _012_
rlabel metal2 s 15410 1768 15410 1768 4 _013_
rlabel metal1 s 16882 4998 16882 4998 4 _014_
rlabel metal2 s 12742 3876 12742 3876 4 _015_
rlabel metal1 s 12512 3366 12512 3366 4 _016_
rlabel metal2 s 2990 3196 2990 3196 4 _017_
rlabel metal1 s 3910 10438 3910 10438 4 _018_
rlabel metal1 s 16977 9010 16977 9010 4 _019_
rlabel metal1 s 15364 12614 15364 12614 4 _020_
rlabel metal1 s 18078 9996 18078 9996 4 _021_
rlabel metal2 s 13202 16677 13202 16677 4 _022_
rlabel metal2 s 17066 7327 17066 7327 4 _023_
rlabel metal1 s 9246 17136 9246 17136 4 _024_
rlabel metal3 s 1587 1020 1587 1020 4 _025_
rlabel metal1 s 3450 8330 3450 8330 4 _026_
rlabel metal1 s 6072 13294 6072 13294 4 _027_
rlabel metal1 s 17894 10676 17894 10676 4 _028_
rlabel metal3 s 14996 6800 14996 6800 4 _029_
rlabel metal2 s 15686 9843 15686 9843 4 _030_
rlabel metal1 s 4646 9520 4646 9520 4 _031_
rlabel metal2 s 5658 7378 5658 7378 4 _032_
rlabel metal2 s 15502 3026 15502 3026 4 _033_
rlabel metal1 s 16560 3026 16560 3026 4 _034_
rlabel metal4 s 16859 3332 16859 3332 4 _035_
rlabel metal1 s 3956 11118 3956 11118 4 _036_
rlabel metal1 s 15226 10778 15226 10778 4 _037_
rlabel metal1 s 18124 11118 18124 11118 4 _038_
rlabel metal1 s 16468 9010 16468 9010 4 _039_
rlabel metal1 s 13938 12954 13938 12954 4 _040_
rlabel metal2 s 17848 12172 17848 12172 4 _041_
rlabel metal1 s 14122 5134 14122 5134 4 _042_
rlabel metal1 s 13294 4114 13294 4114 4 _043_
rlabel metal2 s 5750 6579 5750 6579 4 _044_
rlabel metal1 s 15318 7854 15318 7854 4 _045_
rlabel metal1 s 8050 1598 8050 1598 4 _046_
rlabel metal3 s 11615 14484 11615 14484 4 _047_
rlabel metal4 s 19412 10336 19412 10336 4 _048_
rlabel metal3 s 17526 10013 17526 10013 4 _049_
rlabel metal4 s 18124 7752 18124 7752 4 _050_
rlabel metal1 s 16698 5100 16698 5100 4 _051_
rlabel metal1 s 3910 5202 3910 5202 4 _052_
rlabel metal1 s 14122 7480 14122 7480 4 _053_
rlabel metal2 s 4738 15827 4738 15827 4 _054_
rlabel metal3 s 10028 13668 10028 13668 4 _055_
rlabel metal2 s 11546 7446 11546 7446 4 _056_
rlabel metal2 s 9982 4658 9982 4658 4 _057_
rlabel metal2 s 12466 17068 12466 17068 4 _058_
rlabel metal2 s 10442 16796 10442 16796 4 _059_
rlabel metal1 s 1702 8806 1702 8806 4 _060_
rlabel metal3 s 1219 15300 1219 15300 4 _061_
rlabel metal2 s 1610 8993 1610 8993 4 _062_
rlabel metal1 s 2484 9554 2484 9554 4 _063_
rlabel metal2 s 15318 1751 15318 1751 4 _064_
rlabel metal2 s 16790 17459 16790 17459 4 _065_
rlabel metal2 s 1610 10438 1610 10438 4 _066_
rlabel metal2 s 4186 15708 4186 15708 4 _067_
rlabel metal1 s 14582 3400 14582 3400 4 _068_
rlabel metal2 s 18354 8619 18354 8619 4 _069_
rlabel metal2 s 16606 5831 16606 5831 4 _070_
rlabel metal2 s 7544 9962 7544 9962 4 _071_
rlabel metal2 s 7498 17068 7498 17068 4 _072_
rlabel metal1 s 3128 15334 3128 15334 4 _073_
rlabel metal2 s 18354 15317 18354 15317 4 _074_
rlabel metal1 s 3680 9486 3680 9486 4 _075_
rlabel metal3 s 1932 13396 1932 13396 4 _076_
rlabel metal2 s 4830 2601 4830 2601 4 _077_
rlabel metal2 s 9246 15062 9246 15062 4 _078_
rlabel metal2 s 8970 3910 8970 3910 4 _079_
rlabel metal1 s 10810 12813 10810 12813 4 _080_
rlabel metal1 s 1334 10030 1334 10030 4 _081_
rlabel metal2 s 12466 4624 12466 4624 4 _082_
rlabel metal2 s 6762 12767 6762 12767 4 _083_
rlabel metal1 s 4738 12954 4738 12954 4 _084_
rlabel metal1 s 2070 13158 2070 13158 4 _085_
rlabel metal1 s 11040 16490 11040 16490 4 _086_
rlabel metal2 s 10718 16320 10718 16320 4 _087_
rlabel metal1 s 16514 3468 16514 3468 4 _088_
rlabel metal2 s 15226 4896 15226 4896 4 _089_
rlabel metal2 s 5474 3808 5474 3808 4 _090_
rlabel metal4 s 828 1754 828 1754 4 _091_
rlabel metal2 s 4922 14705 4922 14705 4 _092_
rlabel metal1 s 18768 12206 18768 12206 4 _093_
rlabel metal1 s 17802 12172 17802 12172 4 _094_
rlabel metal2 s 14398 16235 14398 16235 4 _095_
rlabel metal1 s 10350 7310 10350 7310 4 _096_
rlabel metal1 s 10212 7378 10212 7378 4 _097_
rlabel metal1 s 10810 14790 10810 14790 4 _098_
rlabel metal1 s 5014 6324 5014 6324 4 _099_
rlabel metal2 s 5014 4488 5014 4488 4 _100_
rlabel metal2 s 4002 4777 4002 4777 4 _101_
rlabel metal1 s 2254 11866 2254 11866 4 _102_
rlabel metal2 s 14490 16269 14490 16269 4 _103_
rlabel metal1 s 2806 12614 2806 12614 4 _104_
rlabel metal1 s 4416 4658 4416 4658 4 _105_
rlabel metal2 s 13938 15657 13938 15657 4 _106_
rlabel metal1 s 7958 1258 7958 1258 4 _107_
rlabel metal1 s 5198 12852 5198 12852 4 _108_
rlabel metal2 s 2346 1921 2346 1921 4 _109_
rlabel metal2 s 5014 13141 5014 13141 4 _110_
rlabel metal1 s 7268 7854 7268 7854 4 _111_
rlabel metal2 s 16054 2278 16054 2278 4 _112_
rlabel metal1 s 17066 11084 17066 11084 4 _113_
rlabel metal1 s 16698 11152 16698 11152 4 _114_
rlabel metal1 s 13478 12172 13478 12172 4 _115_
rlabel metal2 s 4646 13430 4646 13430 4 _116_
rlabel metal2 s 7682 12682 7682 12682 4 _117_
rlabel metal1 s 12880 12410 12880 12410 4 _118_
rlabel metal1 s 6302 4590 6302 4590 4 _119_
rlabel metal3 s 12834 15453 12834 15453 4 _120_
rlabel metal2 s 2714 3485 2714 3485 4 _121_
rlabel metal3 s 10051 16252 10051 16252 4 _122_
rlabel metal1 s 7038 15674 7038 15674 4 _123_
rlabel metal3 s 11592 16252 11592 16252 4 _124_
rlabel metal3 s 17158 16541 17158 16541 4 _125_
rlabel metal1 s 15870 15878 15870 15878 4 _126_
rlabel metal1 s 14996 7854 14996 7854 4 _127_
rlabel metal1 s 15916 8058 15916 8058 4 _128_
rlabel metal1 s 13018 15028 13018 15028 4 _129_
rlabel metal4 s 8717 2652 8717 2652 4 _130_
rlabel metal2 s 16054 7140 16054 7140 4 _131_
rlabel metal2 s 12650 6817 12650 6817 4 _132_
rlabel metal1 s 17802 5202 17802 5202 4 _133_
rlabel metal1 s 17112 5134 17112 5134 4 _134_
rlabel metal2 s 17526 6052 17526 6052 4 _135_
rlabel metal1 s 13570 6630 13570 6630 4 _136_
rlabel metal2 s 14674 4641 14674 4641 4 _137_
rlabel metal2 s 9062 16762 9062 16762 4 _138_
rlabel metal2 s 9522 16490 9522 16490 4 _139_
rlabel metal1 s 15640 12410 15640 12410 4 _140_
rlabel metal2 s 15410 3247 15410 3247 4 _141_
rlabel metal1 s 4002 12172 4002 12172 4 _142_
rlabel metal2 s 1334 10319 1334 10319 4 _143_
rlabel metal1 s 5198 6902 5198 6902 4 _144_
rlabel metal3 s 7728 14484 7728 14484 4 _145_
rlabel metal1 s 12374 13872 12374 13872 4 _146_
rlabel metal1 s 6256 12342 6256 12342 4 _147_
rlabel metal2 s 12558 9486 12558 9486 4 _148_
rlabel metal1 s 14030 9520 14030 9520 4 _149_
rlabel metal1 s 18078 13260 18078 13260 4 _150_
rlabel metal1 s 14352 14246 14352 14246 4 _151_
rlabel metal2 s 14214 9557 14214 9557 4 _152_
rlabel metal2 s 7038 16031 7038 16031 4 _153_
rlabel metal3 s 5405 15300 5405 15300 4 _154_
rlabel metal1 s 8510 6222 8510 6222 4 _155_
rlabel metal2 s 13754 10302 13754 10302 4 _156_
rlabel metal1 s 6486 14416 6486 14416 4 _157_
rlabel metal1 s 13248 6426 13248 6426 4 _158_
rlabel metal1 s 13110 14348 13110 14348 4 _159_
rlabel metal2 s 8832 14756 8832 14756 4 _160_
rlabel metal1 s 17894 5712 17894 5712 4 _161_
rlabel metal1 s 12880 2278 12880 2278 4 _162_
rlabel metal2 s 12006 2465 12006 2465 4 _163_
rlabel metal1 s 12098 3094 12098 3094 4 _164_
rlabel metal1 s 1886 9588 1886 9588 4 _165_
rlabel metal1 s 1794 9520 1794 9520 4 _166_
rlabel metal2 s 1380 12444 1380 12444 4 _167_
rlabel metal1 s 1426 2414 1426 2414 4 _168_
rlabel metal1 s 2024 2618 2024 2618 4 _169_
rlabel metal1 s 10304 8602 10304 8602 4 _170_
rlabel metal2 s 2576 1428 2576 1428 4 _171_
rlabel metal1 s 7912 9078 7912 9078 4 _172_
rlabel metal2 s 10626 8840 10626 8840 4 _173_
rlabel metal3 s 5405 17068 5405 17068 4 _174_
rlabel metal1 s 2576 5882 2576 5882 4 _175_
rlabel metal2 s 13110 2244 13110 2244 4 _176_
rlabel metal1 s 3680 13294 3680 13294 4 _177_
rlabel metal2 s 13386 14943 13386 14943 4 _178_
rlabel metal2 s 9798 12415 9798 12415 4 _179_
rlabel metal1 s 16100 14586 16100 14586 4 _180_
rlabel metal1 s 6302 11594 6302 11594 4 _181_
rlabel metal3 s 11224 13940 11224 13940 4 _182_
rlabel metal1 s 14398 4590 14398 4590 4 _183_
rlabel metal1 s 6532 8602 6532 8602 4 _184_
rlabel metal1 s 16376 14246 16376 14246 4 _185_
rlabel metal1 s 14904 13294 14904 13294 4 _186_
rlabel metal2 s 14582 4845 14582 4845 4 _187_
rlabel metal1 s 6003 4658 6003 4658 4 _188_
rlabel metal1 s 13570 15674 13570 15674 4 _189_
rlabel metal2 s 2576 12852 2576 12852 4 _190_
rlabel metal1 s 4508 4590 4508 4590 4 _191_
rlabel metal1 s 5382 4794 5382 4794 4 _192_
rlabel metal2 s 3910 13770 3910 13770 4 _193_
rlabel metal3 s 2898 13277 2898 13277 4 _194_
rlabel metal1 s 15226 7786 15226 7786 4 _195_
rlabel metal1 s 2070 4556 2070 4556 4 _196_
rlabel metal1 s 1978 2482 1978 2482 4 _197_
rlabel metal2 s 874 3876 874 3876 4 _198_
rlabel metal1 s 10856 7378 10856 7378 4 _199_
rlabel metal1 s 12650 5304 12650 5304 4 _200_
rlabel metal2 s 17986 2125 17986 2125 4 _201_
rlabel metal2 s 8372 11050 8372 11050 4 _202_
rlabel metal2 s 5934 14076 5934 14076 4 _203_
rlabel metal2 s 1794 16473 1794 16473 4 _204_
rlabel metal1 s 14674 3978 14674 3978 4 _205_
rlabel metal1 s 3864 16218 3864 16218 4 _206_
rlabel metal1 s 1196 12750 1196 12750 4 _207_
rlabel metal1 s 14674 9520 14674 9520 4 _208_
rlabel metal1 s 14858 9554 14858 9554 4 _209_
rlabel metal2 s 6670 5967 6670 5967 4 _210_
rlabel metal1 s 4968 5882 4968 5882 4 _211_
rlabel metal1 s 9200 7854 9200 7854 4 _212_
rlabel metal1 s 3450 13702 3450 13702 4 _213_
rlabel metal4 s 14996 9248 14996 9248 4 _214_
rlabel metal1 s 11684 3910 11684 3910 4 _215_
rlabel metal1 s 3404 6358 3404 6358 4 _216_
rlabel metal2 s 2806 12767 2806 12767 4 _217_
rlabel metal1 s 1978 14450 1978 14450 4 _218_
rlabel metal1 s 13386 11730 13386 11730 4 _219_
rlabel metal2 s 11178 15232 11178 15232 4 _220_
rlabel metal2 s 1978 14161 1978 14161 4 _221_
rlabel metal1 s 13110 11662 13110 11662 4 _222_
rlabel metal2 s 9338 8058 9338 8058 4 _223_
rlabel metal1 s 17710 5270 17710 5270 4 _224_
rlabel metal3 s 15916 12308 15916 12308 4 _225_
rlabel metal2 s 18262 2040 18262 2040 4 _226_
rlabel metal2 s 8050 15674 8050 15674 4 _227_
rlabel metal2 s 9062 7106 9062 7106 4 _228_
rlabel metal1 s 8694 1326 8694 1326 4 _229_
rlabel metal4 s 14628 15288 14628 15288 4 _230_
rlabel metal1 s 11132 2278 11132 2278 4 _231_
rlabel metal1 s 5658 11526 5658 11526 4 _232_
rlabel metal1 s 2254 5576 2254 5576 4 _233_
rlabel metal1 s 1426 5542 1426 5542 4 _234_
rlabel metal2 s 17894 3842 17894 3842 4 _235_
rlabel metal2 s 14214 5593 14214 5593 4 _236_
rlabel metal1 s 6072 2618 6072 2618 4 _237_
rlabel metal1 s 1610 11730 1610 11730 4 _238_
rlabel metal3 s 8878 5253 8878 5253 4 _239_
rlabel metal1 s 7958 3468 7958 3468 4 _240_
rlabel metal1 s 7038 13362 7038 13362 4 _241_
rlabel metal2 s 8234 16830 8234 16830 4 _242_
rlabel metal3 s 13892 1972 13892 1972 4 _243_
rlabel metal1 s 12972 2822 12972 2822 4 _244_
rlabel metal1 s 12918 3162 12918 3162 4 _245_
rlabel metal2 s 15962 18156 15962 18156 4 _246_
rlabel metal2 s 5198 13532 5198 13532 4 _247_
rlabel metal2 s 16882 4369 16882 4369 4 net1
rlabel metal1 s 17158 14960 17158 14960 4 net10
rlabel metal2 s 5198 15844 5198 15844 4 net11
rlabel metal2 s 2254 13192 2254 13192 4 net12
rlabel metal2 s 9798 17374 9798 17374 4 net13
rlabel metal1 s 15226 4624 15226 4624 4 net14
rlabel metal2 s 7406 16660 7406 16660 4 net15
rlabel metal1 s 2070 16626 2070 16626 4 net16
rlabel metal2 s 16882 2142 16882 2142 4 net17
rlabel metal1 s 10764 2482 10764 2482 4 net18
rlabel metal1 s 18124 7854 18124 7854 4 net19
rlabel metal2 s 14030 10574 14030 10574 4 net2
rlabel metal3 s 17342 17187 17342 17187 4 net20
rlabel metal1 s 8004 15334 8004 15334 4 net21
rlabel metal4 s 17940 1564 17940 1564 4 net22
rlabel metal3 s 15870 11237 15870 11237 4 net23
rlabel metal1 s 18262 8908 18262 8908 4 net24
rlabel metal1 s 16054 13430 16054 13430 4 net25
rlabel metal3 s 17917 13940 17917 13940 4 net26
rlabel metal3 s 16813 2516 16813 2516 4 net27
rlabel metal1 s 11178 9146 11178 9146 4 net28
rlabel metal1 s 2162 4114 2162 4114 4 net29
rlabel metal2 s 3266 12903 3266 12903 4 net3
rlabel metal2 s 3634 5406 3634 5406 4 net30
rlabel metal1 s 4922 13294 4922 13294 4 net31
rlabel metal1 s 4370 5678 4370 5678 4 net32
rlabel metal2 s 17526 15453 17526 15453 4 net33
rlabel metal2 s 13570 16456 13570 16456 4 net34
rlabel metal1 s 11224 14382 11224 14382 4 net35
rlabel metal1 s 2162 8500 2162 8500 4 net36
rlabel metal2 s 5198 7276 5198 7276 4 net37
rlabel metal1 s 2300 8806 2300 8806 4 net38
rlabel metal2 s 14306 14433 14306 14433 4 net39
rlabel metal2 s 16698 16252 16698 16252 4 net4
rlabel metal1 s 6992 15538 6992 15538 4 net40
rlabel metal1 s 2806 3434 2806 3434 4 net41
rlabel metal2 s 17434 16711 17434 16711 4 net5
rlabel metal1 s 2024 6834 2024 6834 4 net6
rlabel metal1 s 3128 5202 3128 5202 4 net7
rlabel metal3 s 16238 3672 16238 3672 4 net8
rlabel metal2 s 18170 15283 18170 15283 4 net9
rlabel metal2 s 16606 1588 16606 1588 4 opcode[0]
rlabel metal2 s 9982 1554 9982 1554 4 opcode[1]
rlabel metal2 s 3358 1554 3358 1554 4 opcode[2]
rlabel metal1 s 17710 17306 17710 17306 4 out[0]
rlabel metal2 s 18446 16269 18446 16269 4 out[1]
rlabel metal2 s 18446 13583 18446 13583 4 out[2]
rlabel metal1 s 17204 11254 17204 11254 4 out[3]
rlabel metal3 s 18446 8789 18446 8789 4 out[4]
rlabel metal2 s 18446 6477 18446 6477 4 out[5]
rlabel metal3 s 18446 3893 18446 3893 4 out[6]
rlabel metal3 s 18868 1428 18868 1428 4 out[7]
flabel metal3 s 0 18504 800 18624 0 FreeSans 600 0 0 0 A[0]
port 1 nsew
flabel metal3 s 0 16056 800 16176 0 FreeSans 600 0 0 0 A[1]
port 2 nsew
flabel metal3 s 0 13608 800 13728 0 FreeSans 600 0 0 0 A[2]
port 3 nsew
flabel metal3 s 0 11160 800 11280 0 FreeSans 600 0 0 0 A[3]
port 4 nsew
flabel metal3 s 0 8712 800 8832 0 FreeSans 600 0 0 0 A[4]
port 5 nsew
flabel metal3 s 0 6264 800 6384 0 FreeSans 600 0 0 0 A[5]
port 6 nsew
flabel metal3 s 0 3816 800 3936 0 FreeSans 600 0 0 0 A[6]
port 7 nsew
flabel metal3 s 0 1368 800 1488 0 FreeSans 600 0 0 0 A[7]
port 8 nsew
flabel metal2 s 18602 19200 18658 20000 0 FreeSans 280 90 0 0 B[0]
port 9 nsew
flabel metal2 s 16118 19200 16174 20000 0 FreeSans 280 90 0 0 B[1]
port 10 nsew
flabel metal2 s 13634 19200 13690 20000 0 FreeSans 280 90 0 0 B[2]
port 11 nsew
flabel metal2 s 11150 19200 11206 20000 0 FreeSans 280 90 0 0 B[3]
port 12 nsew
flabel metal2 s 8666 19200 8722 20000 0 FreeSans 280 90 0 0 B[4]
port 13 nsew
flabel metal2 s 6182 19200 6238 20000 0 FreeSans 280 90 0 0 B[5]
port 14 nsew
flabel metal2 s 3698 19200 3754 20000 0 FreeSans 280 90 0 0 B[6]
port 15 nsew
flabel metal2 s 1214 19200 1270 20000 0 FreeSans 280 90 0 0 B[7]
port 16 nsew
flabel metal5 s 1056 13676 18908 13996 0 FreeSans 3200 0 0 0 VGND
port 17 nsew
flabel metal5 s 1056 8676 18908 8996 0 FreeSans 3200 0 0 0 VGND
port 17 nsew
flabel metal5 s 1056 3676 18908 3996 0 FreeSans 3200 0 0 0 VGND
port 17 nsew
flabel metal4 s 17604 2128 17924 17456 0 FreeSans 2400 90 0 0 VGND
port 17 nsew
flabel metal4 s 12604 2128 12924 17456 0 FreeSans 2400 90 0 0 VGND
port 17 nsew
flabel metal4 s 7604 2128 7924 17456 0 FreeSans 2400 90 0 0 VGND
port 17 nsew
flabel metal4 s 2604 2128 2924 17456 0 FreeSans 2400 90 0 0 VGND
port 17 nsew
flabel metal5 s 1056 13016 18908 13336 0 FreeSans 3200 0 0 0 VPWR
port 18 nsew
flabel metal5 s 1056 8016 18908 8336 0 FreeSans 3200 0 0 0 VPWR
port 18 nsew
flabel metal5 s 1056 3016 18908 3336 0 FreeSans 3200 0 0 0 VPWR
port 18 nsew
flabel metal4 s 16944 2128 17264 17456 0 FreeSans 2400 90 0 0 VPWR
port 18 nsew
flabel metal4 s 11944 2128 12264 17456 0 FreeSans 2400 90 0 0 VPWR
port 18 nsew
flabel metal4 s 6944 2128 7264 17456 0 FreeSans 2400 90 0 0 VPWR
port 18 nsew
flabel metal4 s 1944 2128 2264 17456 0 FreeSans 2400 90 0 0 VPWR
port 18 nsew
flabel metal2 s 16578 0 16634 800 0 FreeSans 280 90 0 0 opcode[0]
port 19 nsew
flabel metal2 s 9954 0 10010 800 0 FreeSans 280 90 0 0 opcode[1]
port 20 nsew
flabel metal2 s 3330 0 3386 800 0 FreeSans 280 90 0 0 opcode[2]
port 21 nsew
flabel metal3 s 19200 18504 20000 18624 0 FreeSans 600 0 0 0 out[0]
port 22 nsew
flabel metal3 s 19200 16056 20000 16176 0 FreeSans 600 0 0 0 out[1]
port 23 nsew
flabel metal3 s 19200 13608 20000 13728 0 FreeSans 600 0 0 0 out[2]
port 24 nsew
flabel metal3 s 19200 11160 20000 11280 0 FreeSans 600 0 0 0 out[3]
port 25 nsew
flabel metal3 s 19200 8712 20000 8832 0 FreeSans 600 0 0 0 out[4]
port 26 nsew
flabel metal3 s 19200 6264 20000 6384 0 FreeSans 600 0 0 0 out[5]
port 27 nsew
flabel metal3 s 19200 3816 20000 3936 0 FreeSans 600 0 0 0 out[6]
port 28 nsew
flabel metal3 s 19200 1368 20000 1488 0 FreeSans 600 0 0 0 out[7]
port 29 nsew
<< properties >>
string FIXED_BBOX 0 0 20000 20000
<< end >>
