VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO alu
  CLASS BLOCK ;
  FOREIGN alu ;
  ORIGIN 0.000 0.000 ;
  SIZE 100.000 BY 100.000 ;
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 4.000 93.120 ;
    END
  END A[0]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.280 4.000 80.880 ;
    END
  END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 4.000 56.400 ;
    END
  END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 4.000 44.160 ;
    END
  END A[4]
  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 4.000 31.920 ;
    END
  END A[5]
  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 4.000 19.680 ;
    END
  END A[6]
  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END A[7]
  PIN B[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 93.010 96.000 93.290 100.000 ;
    END
  END B[0]
  PIN B[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 80.590 96.000 80.870 100.000 ;
    END
  END B[1]
  PIN B[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 68.170 96.000 68.450 100.000 ;
    END
  END B[2]
  PIN B[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 55.750 96.000 56.030 100.000 ;
    END
  END B[3]
  PIN B[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 43.330 96.000 43.610 100.000 ;
    END
  END B[4]
  PIN B[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 30.910 96.000 31.190 100.000 ;
    END
  END B[5]
  PIN B[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 18.490 96.000 18.770 100.000 ;
    END
  END B[6]
  PIN B[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 6.070 96.000 6.350 100.000 ;
    END
  END B[7]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 13.020 10.640 14.620 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 38.020 10.640 39.620 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 63.020 10.640 64.620 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 88.020 10.640 89.620 87.280 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 18.380 94.540 19.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 43.380 94.540 44.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 68.380 94.540 69.980 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 9.720 10.640 11.320 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 34.720 10.640 36.320 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 59.720 10.640 61.320 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 84.720 10.640 86.320 87.280 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 15.080 94.540 16.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 40.080 94.540 41.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 65.080 94.540 66.680 ;
    END
  END VPWR
  PIN opcode[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 82.890 0.000 83.170 4.000 ;
    END
  END opcode[0]
  PIN opcode[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 4.000 ;
    END
  END opcode[1]
  PIN opcode[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 16.650 0.000 16.930 4.000 ;
    END
  END opcode[2]
  PIN out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 96.000 92.520 100.000 93.120 ;
    END
  END out[0]
  PIN out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 96.000 80.280 100.000 80.880 ;
    END
  END out[1]
  PIN out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 96.000 68.040 100.000 68.640 ;
    END
  END out[2]
  PIN out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 96.000 55.800 100.000 56.400 ;
    END
  END out[3]
  PIN out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 96.000 43.560 100.000 44.160 ;
    END
  END out[4]
  PIN out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 96.000 31.320 100.000 31.920 ;
    END
  END out[5]
  PIN out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 96.000 19.080 100.000 19.680 ;
    END
  END out[6]
  PIN out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 96.000 6.840 100.000 7.440 ;
    END
  END out[7]
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 94.490 87.125 ;
      LAYER li1 ;
        RECT 5.520 10.795 94.300 87.125 ;
      LAYER met1 ;
        RECT 0.530 2.420 97.910 94.140 ;
      LAYER met2 ;
        RECT 0.550 95.720 5.790 96.000 ;
        RECT 6.630 95.720 18.210 96.000 ;
        RECT 19.050 95.720 30.630 96.000 ;
        RECT 31.470 95.720 43.050 96.000 ;
        RECT 43.890 95.720 55.470 96.000 ;
        RECT 56.310 95.720 67.890 96.000 ;
        RECT 68.730 95.720 80.310 96.000 ;
        RECT 81.150 95.720 92.730 96.000 ;
        RECT 93.570 95.720 97.880 96.000 ;
        RECT 0.550 4.280 97.880 95.720 ;
        RECT 0.550 2.195 16.370 4.280 ;
        RECT 17.210 2.195 49.490 4.280 ;
        RECT 50.330 2.195 82.610 4.280 ;
        RECT 83.450 2.195 97.880 4.280 ;
      LAYER met3 ;
        RECT 0.525 93.520 97.250 93.665 ;
        RECT 4.400 92.120 95.600 93.520 ;
        RECT 0.525 81.280 97.250 92.120 ;
        RECT 4.400 79.880 95.600 81.280 ;
        RECT 0.525 69.040 97.250 79.880 ;
        RECT 4.400 67.640 95.600 69.040 ;
        RECT 0.525 56.800 97.250 67.640 ;
        RECT 4.400 55.400 95.600 56.800 ;
        RECT 0.525 44.560 97.250 55.400 ;
        RECT 4.400 43.160 95.600 44.560 ;
        RECT 0.525 32.320 97.250 43.160 ;
        RECT 4.400 30.920 95.600 32.320 ;
        RECT 0.525 20.080 97.250 30.920 ;
        RECT 4.400 18.680 95.600 20.080 ;
        RECT 0.525 7.840 97.250 18.680 ;
        RECT 4.400 6.440 95.600 7.840 ;
        RECT 0.525 2.215 97.250 6.440 ;
      LAYER met4 ;
        RECT 3.975 87.680 97.650 93.665 ;
        RECT 3.975 10.240 9.320 87.680 ;
        RECT 11.720 10.240 12.620 87.680 ;
        RECT 15.020 10.240 34.320 87.680 ;
        RECT 36.720 10.240 37.620 87.680 ;
        RECT 40.020 10.240 59.320 87.680 ;
        RECT 61.720 10.240 62.620 87.680 ;
        RECT 65.020 10.240 84.320 87.680 ;
        RECT 86.720 10.240 87.620 87.680 ;
        RECT 90.020 10.240 97.650 87.680 ;
        RECT 3.975 2.215 97.650 10.240 ;
      LAYER met5 ;
        RECT 4.260 71.580 97.860 84.100 ;
        RECT 96.140 63.480 97.860 71.580 ;
        RECT 4.260 46.580 97.860 63.480 ;
        RECT 96.140 38.480 97.860 46.580 ;
        RECT 4.260 21.580 97.860 38.480 ;
        RECT 96.140 13.480 97.860 21.580 ;
        RECT 4.260 4.300 97.860 13.480 ;
  END
END alu
END LIBRARY

