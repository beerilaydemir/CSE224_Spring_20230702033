* NGSPICE file created from ZeroToFiveCounter.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

.subckt ZeroToFiveCounter AN[0] AN[1] AN[2] AN[3] AN[4] AN[5] AN[6] AN[7] VGND VPWR
+ clk count[0] count[1] count[2] count[3] rst
X_363_ clknet_2_2__leaf_clk _026_ _040_ VGND VGND VPWR VPWR one_second_counter\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_294_ _148_ one_second_counter\[20\] _150_ VGND VGND VPWR VPWR _152_ sky130_fd_sc_hd__nand3_1
XFILLER_0_13_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_0_Left_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_346_ _169_ VGND VGND VPWR VPWR _054_ sky130_fd_sc_hd__inv_2
X_277_ one_second_counter\[16\] _135_ VGND VGND VPWR VPWR _139_ sky130_fd_sc_hd__or2_1
X_200_ net17 VGND VGND VPWR VPWR _078_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_329_ _168_ VGND VGND VPWR VPWR _038_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_95 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_293_ _148_ _150_ _151_ _086_ VGND VGND VPWR VPWR _010_ sky130_fd_sc_hd__o211a_1
X_362_ clknet_2_2__leaf_clk _025_ _039_ VGND VGND VPWR VPWR one_second_counter\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_276_ one_second_counter\[16\] _135_ VGND VGND VPWR VPWR _138_ sky130_fd_sc_hd__nand2_1
X_345_ _169_ VGND VGND VPWR VPWR _053_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_259_ one_second_counter\[12\] one_second_counter\[11\] _121_ VGND VGND VPWR VPWR
+ _125_ sky130_fd_sc_hd__and3_1
X_328_ _168_ VGND VGND VPWR VPWR _037_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_292_ _148_ _150_ VGND VGND VPWR VPWR _151_ sky130_fd_sc_hd__nand2_1
X_361_ clknet_2_0__leaf_clk _024_ _038_ VGND VGND VPWR VPWR one_second_counter\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_275_ _137_ VGND VGND VPWR VPWR _006_ sky130_fd_sc_hd__clkbuf_1
X_344_ _169_ VGND VGND VPWR VPWR _052_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_258_ one_second_counter\[12\] _122_ VGND VGND VPWR VPWR _124_ sky130_fd_sc_hd__or2_1
X_189_ net3 net2 _068_ net4 VGND VGND VPWR VPWR _070_ sky130_fd_sc_hd__a31o_1
X_327_ net1 VGND VGND VPWR VPWR _168_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_5_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_16_Left_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_64 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_291_ _149_ VGND VGND VPWR VPWR _150_ sky130_fd_sc_hd__buf_2
XFILLER_0_7_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_360_ clknet_2_0__leaf_clk _023_ _037_ VGND VGND VPWR VPWR one_second_counter\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_19_Left_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_274_ _096_ _133_ _136_ VGND VGND VPWR VPWR _137_ sky130_fd_sc_hd__and3_1
X_343_ _169_ VGND VGND VPWR VPWR _051_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_4_Left_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_188_ net14 _069_ VGND VGND VPWR VPWR _061_ sky130_fd_sc_hd__xor2_1
X_326_ _167_ VGND VGND VPWR VPWR _036_ sky130_fd_sc_hd__inv_2
X_257_ net18 _120_ _123_ _086_ VGND VGND VPWR VPWR _002_ sky130_fd_sc_hd__o211a_1
XFILLER_0_19_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_309_ _079_ _159_ _146_ _162_ _086_ VGND VGND VPWR VPWR _016_ sky130_fd_sc_hd__o311a_1
XPHY_EDGE_ROW_7_Left_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_15_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_290_ one_second_counter\[11\] _134_ _121_ _145_ VGND VGND VPWR VPWR _149_ sky130_fd_sc_hd__and4_1
X_342_ _169_ VGND VGND VPWR VPWR _050_ sky130_fd_sc_hd__inv_2
X_273_ _135_ VGND VGND VPWR VPWR _136_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_20_Left_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_187_ net4 net3 net2 _068_ VGND VGND VPWR VPWR _069_ sky130_fd_sc_hd__and4_1
X_325_ _167_ VGND VGND VPWR VPWR _035_ sky130_fd_sc_hd__inv_2
X_256_ _122_ VGND VGND VPWR VPWR _123_ sky130_fd_sc_hd__inv_2
Xclkload0 clknet_2_0__leaf_clk VGND VGND VPWR VPWR clkload0/X sky130_fd_sc_hd__clkbuf_4
X_308_ _148_ _173_ _150_ one_second_counter\[24\] VGND VGND VPWR VPWR _162_ sky130_fd_sc_hd__a31o_1
X_239_ _108_ VGND VGND VPWR VPWR _109_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_272_ one_second_counter\[11\] _134_ _121_ VGND VGND VPWR VPWR _135_ sky130_fd_sc_hd__and3_2
X_341_ _169_ VGND VGND VPWR VPWR _049_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_324_ _167_ VGND VGND VPWR VPWR _034_ sky130_fd_sc_hd__inv_2
X_186_ _172_ _063_ _065_ _067_ VGND VGND VPWR VPWR _068_ sky130_fd_sc_hd__and4_1
X_255_ one_second_counter\[11\] _121_ VGND VGND VPWR VPWR _122_ sky130_fd_sc_hd__and2_1
Xclkload1 clknet_2_2__leaf_clk VGND VGND VPWR VPWR clkload1/X sky130_fd_sc_hd__clkbuf_4
X_238_ one_second_counter\[8\] _170_ _171_ VGND VGND VPWR VPWR _108_ sky130_fd_sc_hd__and3_1
X_307_ _159_ _146_ _161_ _086_ VGND VGND VPWR VPWR _015_ sky130_fd_sc_hd__o211a_1
XFILLER_0_15_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_6_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_340_ _169_ VGND VGND VPWR VPWR _048_ sky130_fd_sc_hd__inv_2
X_271_ one_second_counter\[12\] _062_ VGND VGND VPWR VPWR _134_ sky130_fd_sc_hd__and2_1
X_323_ _167_ VGND VGND VPWR VPWR _033_ sky130_fd_sc_hd__inv_2
X_185_ one_second_counter\[12\] _066_ VGND VGND VPWR VPWR _067_ sky130_fd_sc_hd__nor2_1
X_254_ one_second_counter\[8\] _170_ _171_ _116_ VGND VGND VPWR VPWR _121_ sky130_fd_sc_hd__and4_1
Xclkload2 clknet_2_3__leaf_clk VGND VGND VPWR VPWR clkload2/X sky130_fd_sc_hd__clkbuf_4
X_237_ _107_ VGND VGND VPWR VPWR _024_ sky130_fd_sc_hd__clkbuf_1
X_306_ _148_ _160_ _150_ net16 VGND VGND VPWR VPWR _161_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_6_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_270_ one_second_counter\[13\] one_second_counter\[14\] _125_ one_second_counter\[15\]
+ VGND VGND VPWR VPWR _133_ sky130_fd_sc_hd__a31o_1
XFILLER_0_4_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_322_ _167_ VGND VGND VPWR VPWR _032_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_184_ one_second_counter\[8\] one_second_counter\[9\] one_second_counter\[10\] one_second_counter\[11\]
+ VGND VGND VPWR VPWR _066_ sky130_fd_sc_hd__or4_1
X_253_ one_second_counter\[9\] one_second_counter\[10\] _108_ VGND VGND VPWR VPWR
+ _120_ sky130_fd_sc_hd__and3_1
X_236_ _172_ _085_ _106_ VGND VGND VPWR VPWR _107_ sky130_fd_sc_hd__and3b_1
X_305_ one_second_counter\[20\] one_second_counter\[21\] one_second_counter\[22\]
+ VGND VGND VPWR VPWR _160_ sky130_fd_sc_hd__and3_1
X_219_ one_second_counter\[0\] one_second_counter\[1\] one_second_counter\[2\] one_second_counter\[3\]
+ VGND VGND VPWR VPWR _094_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_11_Left_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_321_ _167_ VGND VGND VPWR VPWR _031_ sky130_fd_sc_hd__inv_2
X_183_ one_second_counter\[25\] _064_ VGND VGND VPWR VPWR _065_ sky130_fd_sc_hd__nor2_1
X_252_ _119_ VGND VGND VPWR VPWR _001_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_235_ one_second_counter\[5\] one_second_counter\[6\] _097_ one_second_counter\[7\]
+ VGND VGND VPWR VPWR _106_ sky130_fd_sc_hd__a31o_1
X_304_ _148_ _173_ VGND VGND VPWR VPWR _159_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_218_ _093_ VGND VGND VPWR VPWR _019_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_2_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_4_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_320_ _167_ VGND VGND VPWR VPWR _030_ sky130_fd_sc_hd__inv_2
X_182_ one_second_counter\[26\] one_second_counter\[24\] VGND VGND VPWR VPWR _064_
+ sky130_fd_sc_hd__nand2_1
X_251_ _096_ _117_ _118_ VGND VGND VPWR VPWR _119_ sky130_fd_sc_hd__and3_1
X_303_ _157_ _151_ _158_ _086_ VGND VGND VPWR VPWR _014_ sky130_fd_sc_hd__o211a_1
X_234_ _104_ _098_ _105_ _086_ VGND VGND VPWR VPWR _023_ sky130_fd_sc_hd__o211a_1
XFILLER_0_21_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_217_ _091_ _085_ _092_ VGND VGND VPWR VPWR _093_ sky130_fd_sc_hd__and3_1
XFILLER_0_22_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_250_ one_second_counter\[10\] _112_ VGND VGND VPWR VPWR _118_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_181_ _173_ _174_ _062_ VGND VGND VPWR VPWR _063_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_13_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_379_ clknet_2_1__leaf_clk _017_ _056_ VGND VGND VPWR VPWR one_second_counter\[25\]
+ sky130_fd_sc_hd__dfrtp_2
X_233_ one_second_counter\[4\] one_second_counter\[5\] _170_ one_second_counter\[6\]
+ VGND VGND VPWR VPWR _105_ sky130_fd_sc_hd__a31o_1
X_302_ _148_ one_second_counter\[20\] one_second_counter\[21\] _150_ one_second_counter\[22\]
+ VGND VGND VPWR VPWR _158_ sky130_fd_sc_hd__a41o_1
X_216_ one_second_counter\[0\] one_second_counter\[1\] one_second_counter\[2\] VGND
+ VGND VPWR VPWR _092_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_15_Left_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_94 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_180_ one_second_counter\[13\] one_second_counter\[14\] one_second_counter\[15\]
+ VGND VGND VPWR VPWR _062_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_18_Left_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_378_ clknet_2_1__leaf_clk _016_ _055_ VGND VGND VPWR VPWR one_second_counter\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_3_Left_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_301_ one_second_counter\[20\] one_second_counter\[21\] one_second_counter\[22\]
+ VGND VGND VPWR VPWR _157_ sky130_fd_sc_hd__nand3_1
XFILLER_0_5_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_232_ one_second_counter\[5\] one_second_counter\[6\] VGND VGND VPWR VPWR _104_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_215_ one_second_counter\[0\] one_second_counter\[1\] one_second_counter\[2\] VGND
+ VGND VPWR VPWR _091_ sky130_fd_sc_hd__nand3_1
XFILLER_0_12_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_377_ clknet_2_3__leaf_clk _015_ _054_ VGND VGND VPWR VPWR one_second_counter\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_300_ _155_ _151_ _156_ _086_ VGND VGND VPWR VPWR _013_ sky130_fd_sc_hd__o211a_1
X_231_ _103_ VGND VGND VPWR VPWR _022_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput1 rst VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_1
XFILLER_0_20_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_214_ _090_ VGND VGND VPWR VPWR _011_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_376_ clknet_2_3__leaf_clk _014_ _053_ VGND VGND VPWR VPWR one_second_counter\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_230_ _096_ _101_ _102_ VGND VGND VPWR VPWR _103_ sky130_fd_sc_hd__and3_1
X_359_ clknet_2_0__leaf_clk _022_ _036_ VGND VGND VPWR VPWR one_second_counter\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_19_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_213_ _088_ _085_ _089_ VGND VGND VPWR VPWR _090_ sky130_fd_sc_hd__and3_1
XFILLER_0_22_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_375_ clknet_2_3__leaf_clk _013_ _052_ VGND VGND VPWR VPWR one_second_counter\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_358_ clknet_2_0__leaf_clk _021_ _035_ VGND VGND VPWR VPWR one_second_counter\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_289_ one_second_counter\[19\] VGND VGND VPWR VPWR _148_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_10_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_212_ one_second_counter\[0\] one_second_counter\[1\] VGND VGND VPWR VPWR _089_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_374_ clknet_2_1__leaf_clk _012_ _051_ VGND VGND VPWR VPWR one_second_counter\[20\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_18_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_357_ clknet_2_0__leaf_clk _020_ _034_ VGND VGND VPWR VPWR one_second_counter\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_2_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_10_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_288_ _147_ VGND VGND VPWR VPWR _009_ sky130_fd_sc_hd__clkbuf_1
X_211_ one_second_counter\[0\] one_second_counter\[1\] VGND VGND VPWR VPWR _088_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_10_Left_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_373_ clknet_2_3__leaf_clk _010_ _050_ VGND VGND VPWR VPWR one_second_counter\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_356_ clknet_2_0__leaf_clk _019_ _033_ VGND VGND VPWR VPWR one_second_counter\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_287_ _085_ _144_ _146_ VGND VGND VPWR VPWR _147_ sky130_fd_sc_hd__and3_1
XFILLER_0_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_210_ _087_ VGND VGND VPWR VPWR _000_ sky130_fd_sc_hd__clkbuf_1
X_339_ _169_ VGND VGND VPWR VPWR _047_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_372_ clknet_2_3__leaf_clk _009_ _049_ VGND VGND VPWR VPWR one_second_counter\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_355_ clknet_2_0__leaf_clk _011_ _032_ VGND VGND VPWR VPWR one_second_counter\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_1_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_286_ _135_ _145_ VGND VGND VPWR VPWR _146_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_269_ _131_ _126_ _132_ _086_ VGND VGND VPWR VPWR _005_ sky130_fd_sc_hd__o211a_1
X_338_ net1 VGND VGND VPWR VPWR _169_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_11_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_371_ clknet_2_3__leaf_clk _008_ _048_ VGND VGND VPWR VPWR one_second_counter\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_285_ one_second_counter\[17\] one_second_counter\[16\] one_second_counter\[18\]
+ VGND VGND VPWR VPWR _145_ sky130_fd_sc_hd__and3_1
XFILLER_0_1_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_354_ clknet_2_0__leaf_clk _000_ _031_ VGND VGND VPWR VPWR one_second_counter\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_1_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_337_ _168_ VGND VGND VPWR VPWR _046_ sky130_fd_sc_hd__inv_2
X_268_ one_second_counter\[13\] _125_ one_second_counter\[14\] VGND VGND VPWR VPWR
+ _132_ sky130_fd_sc_hd__a21o_1
X_199_ _077_ VGND VGND VPWR VPWR _058_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_14_Left_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_370_ clknet_2_3__leaf_clk _007_ _047_ VGND VGND VPWR VPWR one_second_counter\[16\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_17_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_17_Left_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_284_ one_second_counter\[17\] one_second_counter\[16\] _135_ one_second_counter\[18\]
+ VGND VGND VPWR VPWR _144_ sky130_fd_sc_hd__a31o_1
X_353_ clknet_2_1__leaf_clk _061_ _030_ VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_2_Left_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_336_ _168_ VGND VGND VPWR VPWR _045_ sky130_fd_sc_hd__inv_2
X_267_ one_second_counter\[13\] one_second_counter\[14\] VGND VGND VPWR VPWR _131_
+ sky130_fd_sc_hd__nand2_1
X_198_ _075_ _071_ _076_ VGND VGND VPWR VPWR _077_ sky130_fd_sc_hd__and3_1
X_319_ _167_ VGND VGND VPWR VPWR _029_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_7_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_283_ _143_ VGND VGND VPWR VPWR _008_ sky130_fd_sc_hd__clkbuf_1
X_352_ clknet_2_1__leaf_clk _060_ _029_ VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_335_ _168_ VGND VGND VPWR VPWR _044_ sky130_fd_sc_hd__inv_2
X_266_ _130_ VGND VGND VPWR VPWR _004_ sky130_fd_sc_hd__clkbuf_1
X_197_ net2 _068_ VGND VGND VPWR VPWR _076_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_112 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_318_ _167_ VGND VGND VPWR VPWR _028_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_7_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_249_ _108_ _116_ VGND VGND VPWR VPWR _117_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_22_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1 net5 VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_282_ _096_ _141_ _142_ VGND VGND VPWR VPWR _143_ sky130_fd_sc_hd__and3_1
X_351_ clknet_2_1__leaf_clk _059_ _028_ VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_334_ _168_ VGND VGND VPWR VPWR _043_ sky130_fd_sc_hd__inv_2
X_265_ _096_ _128_ _129_ VGND VGND VPWR VPWR _130_ sky130_fd_sc_hd__and3_1
X_196_ net15 _075_ VGND VGND VPWR VPWR _059_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_179_ one_second_counter\[17\] one_second_counter\[19\] one_second_counter\[18\]
+ one_second_counter\[16\] VGND VGND VPWR VPWR _174_ sky130_fd_sc_hd__and4bb_1
X_317_ _167_ VGND VGND VPWR VPWR _027_ sky130_fd_sc_hd__inv_2
X_248_ one_second_counter\[9\] one_second_counter\[10\] VGND VGND VPWR VPWR _116_
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_22_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_2_2__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_19_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2 net3 VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_281_ one_second_counter\[16\] _135_ one_second_counter\[17\] VGND VGND VPWR VPWR
+ _142_ sky130_fd_sc_hd__a21o_1
X_350_ clknet_2_1__leaf_clk _058_ _027_ VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_264_ one_second_counter\[13\] _125_ VGND VGND VPWR VPWR _129_ sky130_fd_sc_hd__nand2_1
X_195_ one_second_counter\[25\] _064_ _074_ net2 VGND VGND VPWR VPWR _075_ sky130_fd_sc_hd__or4b_1
X_333_ _168_ VGND VGND VPWR VPWR _042_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_6_Left_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_247_ _115_ VGND VGND VPWR VPWR _026_ sky130_fd_sc_hd__clkbuf_1
X_316_ net1 VGND VGND VPWR VPWR _167_ sky130_fd_sc_hd__buf_4
X_178_ one_second_counter\[20\] one_second_counter\[21\] one_second_counter\[22\]
+ one_second_counter\[23\] VGND VGND VPWR VPWR _173_ sky130_fd_sc_hd__and4_1
XFILLER_0_18_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_9_Left_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold3 one_second_counter\[23\] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__dlygate4sd3_1
X_280_ one_second_counter\[17\] one_second_counter\[16\] _135_ VGND VGND VPWR VPWR
+ _141_ sky130_fd_sc_hd__nand3_1
XFILLER_0_22_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_22_Left_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_263_ one_second_counter\[13\] _125_ VGND VGND VPWR VPWR _128_ sky130_fd_sc_hd__or2_1
X_194_ _172_ _173_ _174_ _073_ VGND VGND VPWR VPWR _074_ sky130_fd_sc_hd__nand4_1
X_332_ _168_ VGND VGND VPWR VPWR _041_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_246_ _096_ _113_ _114_ VGND VGND VPWR VPWR _115_ sky130_fd_sc_hd__and3_1
X_315_ _078_ _165_ _086_ VGND VGND VPWR VPWR _018_ sky130_fd_sc_hd__a21boi_1
X_177_ _170_ _171_ VGND VGND VPWR VPWR _172_ sky130_fd_sc_hd__and2_1
X_229_ one_second_counter\[5\] _097_ VGND VGND VPWR VPWR _102_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4 one_second_counter\[26\] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_331_ _168_ VGND VGND VPWR VPWR _040_ sky130_fd_sc_hd__inv_2
X_262_ _127_ VGND VGND VPWR VPWR _003_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_60 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_193_ _066_ one_second_counter\[12\] _062_ VGND VGND VPWR VPWR _073_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_2_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_314_ _166_ VGND VGND VPWR VPWR _017_ sky130_fd_sc_hd__clkbuf_1
X_176_ one_second_counter\[4\] one_second_counter\[5\] one_second_counter\[6\] one_second_counter\[7\]
+ VGND VGND VPWR VPWR _171_ sky130_fd_sc_hd__and4_1
X_245_ one_second_counter\[9\] _108_ VGND VGND VPWR VPWR _114_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_228_ one_second_counter\[5\] _097_ VGND VGND VPWR VPWR _101_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_4_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5 one_second_counter\[11\] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_261_ _096_ _124_ _126_ VGND VGND VPWR VPWR _127_ sky130_fd_sc_hd__and3_1
X_192_ _072_ VGND VGND VPWR VPWR _060_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_330_ _168_ VGND VGND VPWR VPWR _039_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_244_ _112_ VGND VGND VPWR VPWR _113_ sky130_fd_sc_hd__inv_2
X_175_ one_second_counter\[0\] one_second_counter\[1\] one_second_counter\[2\] one_second_counter\[3\]
+ VGND VGND VPWR VPWR _170_ sky130_fd_sc_hd__and4_2
X_313_ _085_ _163_ _165_ VGND VGND VPWR VPWR _166_ sky130_fd_sc_hd__and3_1
XFILLER_0_3_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_227_ _100_ VGND VGND VPWR VPWR _021_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_260_ _125_ VGND VGND VPWR VPWR _126_ sky130_fd_sc_hd__inv_2
X_191_ _069_ _070_ _071_ VGND VGND VPWR VPWR _072_ sky130_fd_sc_hd__and3b_1
XFILLER_0_6_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_312_ _079_ _164_ _159_ _150_ VGND VGND VPWR VPWR _165_ sky130_fd_sc_hd__or4b_1
X_243_ one_second_counter\[9\] _108_ VGND VGND VPWR VPWR _112_ sky130_fd_sc_hd__and2_1
X_226_ _096_ _098_ _099_ VGND VGND VPWR VPWR _100_ sky130_fd_sc_hd__and3_1
X_209_ one_second_counter\[0\] _086_ VGND VGND VPWR VPWR _087_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_13_Left_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_190_ net5 net3 net2 net4 VGND VGND VPWR VPWR _071_ sky130_fd_sc_hd__or4b_1
XFILLER_0_12_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_1_Left_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_311_ one_second_counter\[25\] VGND VGND VPWR VPWR _164_ sky130_fd_sc_hd__inv_2
X_242_ _111_ VGND VGND VPWR VPWR _025_ sky130_fd_sc_hd__clkbuf_1
X_225_ one_second_counter\[4\] _170_ VGND VGND VPWR VPWR _099_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_208_ _085_ VGND VGND VPWR VPWR _086_ sky130_fd_sc_hd__buf_2
XFILLER_0_0_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_2_3__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_310_ _148_ one_second_counter\[24\] _173_ _150_ one_second_counter\[25\] VGND VGND
+ VPWR VPWR _163_ sky130_fd_sc_hd__a41o_1
X_241_ _096_ _109_ _110_ VGND VGND VPWR VPWR _111_ sky130_fd_sc_hd__and3_1
XFILLER_0_3_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_224_ _097_ VGND VGND VPWR VPWR _098_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_207_ _078_ _079_ _083_ _084_ VGND VGND VPWR VPWR _085_ sky130_fd_sc_hd__o31a_2
XFILLER_0_0_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_116 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XZeroToFiveCounter_10 VGND VGND VPWR VPWR AN[1] ZeroToFiveCounter_10/LO sky130_fd_sc_hd__conb_1
X_240_ one_second_counter\[8\] _172_ VGND VGND VPWR VPWR _110_ sky130_fd_sc_hd__or2_1
X_369_ clknet_2_2__leaf_clk _006_ _046_ VGND VGND VPWR VPWR one_second_counter\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_223_ one_second_counter\[4\] _170_ VGND VGND VPWR VPWR _097_ sky130_fd_sc_hd__and2_1
X_206_ one_second_counter\[26\] one_second_counter\[25\] VGND VGND VPWR VPWR _084_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XZeroToFiveCounter_11 VGND VGND VPWR VPWR AN[2] ZeroToFiveCounter_11/LO sky130_fd_sc_hd__conb_1
XFILLER_0_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_368_ clknet_2_2__leaf_clk _005_ _045_ VGND VGND VPWR VPWR one_second_counter\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_299_ _148_ one_second_counter\[20\] _150_ one_second_counter\[21\] VGND VGND VPWR
+ VPWR _156_ sky130_fd_sc_hd__a31o_1
XFILLER_0_2_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_5_Left_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_222_ _085_ VGND VGND VPWR VPWR _096_ sky130_fd_sc_hd__clkbuf_2
X_205_ _063_ _080_ _082_ VGND VGND VPWR VPWR _083_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Left_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XZeroToFiveCounter_6 VGND VGND VPWR VPWR ZeroToFiveCounter_6/HI AN[0] sky130_fd_sc_hd__conb_1
XFILLER_0_6_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XZeroToFiveCounter_12 VGND VGND VPWR VPWR AN[6] ZeroToFiveCounter_12/LO sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_2_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput2 net2 VGND VGND VPWR VPWR count[0] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_21_Left_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_367_ clknet_2_2__leaf_clk _004_ _044_ VGND VGND VPWR VPWR one_second_counter\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_298_ one_second_counter\[20\] one_second_counter\[21\] VGND VGND VPWR VPWR _155_
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_12_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_221_ _095_ VGND VGND VPWR VPWR _020_ sky130_fd_sc_hd__clkbuf_1
X_204_ _173_ _081_ VGND VGND VPWR VPWR _082_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XZeroToFiveCounter_7 VGND VGND VPWR VPWR ZeroToFiveCounter_7/HI AN[3] sky130_fd_sc_hd__conb_1
XFILLER_0_6_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XZeroToFiveCounter_13 VGND VGND VPWR VPWR AN[7] ZeroToFiveCounter_13/LO sky130_fd_sc_hd__conb_1
Xoutput3 net3 VGND VGND VPWR VPWR count[1] sky130_fd_sc_hd__buf_2
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_366_ clknet_2_2__leaf_clk _003_ _043_ VGND VGND VPWR VPWR one_second_counter\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_297_ _154_ VGND VGND VPWR VPWR _012_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_59 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_220_ _170_ _085_ _094_ VGND VGND VPWR VPWR _095_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_12_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_349_ net1 VGND VGND VPWR VPWR _057_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_203_ one_second_counter\[17\] one_second_counter\[18\] one_second_counter\[19\]
+ VGND VGND VPWR VPWR _081_ sky130_fd_sc_hd__a21o_1
XFILLER_0_19_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XZeroToFiveCounter_8 VGND VGND VPWR VPWR ZeroToFiveCounter_8/HI AN[4] sky130_fd_sc_hd__conb_1
XFILLER_0_13_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput4 net4 VGND VGND VPWR VPWR count[2] sky130_fd_sc_hd__buf_2
XFILLER_0_5_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_296_ _085_ _152_ _153_ VGND VGND VPWR VPWR _154_ sky130_fd_sc_hd__and3_1
X_365_ clknet_2_2__leaf_clk _002_ _042_ VGND VGND VPWR VPWR one_second_counter\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_279_ _140_ VGND VGND VPWR VPWR _007_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_348_ _169_ VGND VGND VPWR VPWR _056_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_202_ _170_ _171_ _066_ one_second_counter\[12\] VGND VGND VPWR VPWR _080_ sky130_fd_sc_hd__a211o_1
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_50 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XZeroToFiveCounter_9 VGND VGND VPWR VPWR ZeroToFiveCounter_9/HI AN[5] sky130_fd_sc_hd__conb_1
XFILLER_0_21_60 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput5 net5 VGND VGND VPWR VPWR count[3] sky130_fd_sc_hd__buf_2
XFILLER_0_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_295_ _148_ _150_ one_second_counter\[20\] VGND VGND VPWR VPWR _153_ sky130_fd_sc_hd__a21o_1
X_364_ clknet_2_2__leaf_clk _001_ _041_ VGND VGND VPWR VPWR one_second_counter\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_94 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_278_ _096_ _138_ _139_ VGND VGND VPWR VPWR _140_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_347_ _169_ VGND VGND VPWR VPWR _055_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_201_ one_second_counter\[24\] VGND VGND VPWR VPWR _079_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_62 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_18_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_12_Left_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_380_ clknet_2_1__leaf_clk _018_ _057_ VGND VGND VPWR VPWR one_second_counter\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
.ends

