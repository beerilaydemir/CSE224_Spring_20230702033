magic
tech sky130A
magscale 1 2
timestamp 1747771759
<< checkpaint >>
rect -3932 -3932 18819 18668
<< viali >>
rect 5733 13889 5767 13923
rect 6561 13889 6595 13923
rect 1409 13821 1443 13855
rect 5825 13821 5859 13855
rect 5917 13821 5951 13855
rect 6009 13821 6043 13855
rect 9505 13821 9539 13855
rect 9781 13821 9815 13855
rect 13369 13821 13403 13855
rect 6193 13685 6227 13719
rect 6377 13685 6411 13719
rect 8033 13685 8067 13719
rect 3985 13481 4019 13515
rect 4261 13481 4295 13515
rect 6837 13481 6871 13515
rect 7389 13481 7423 13515
rect 7849 13481 7883 13515
rect 9045 13481 9079 13515
rect 9413 13481 9447 13515
rect 9597 13481 9631 13515
rect 7573 13413 7607 13447
rect 8033 13413 8067 13447
rect 5089 13345 5123 13379
rect 5365 13345 5399 13379
rect 3341 13277 3375 13311
rect 3433 13277 3467 13311
rect 4445 13277 4479 13311
rect 4813 13277 4847 13311
rect 4997 13277 5031 13311
rect 7113 13277 7147 13311
rect 8125 13277 8159 13311
rect 8309 13277 8343 13311
rect 8769 13277 8803 13311
rect 8953 13277 8987 13311
rect 9137 13277 9171 13311
rect 9229 13277 9263 13311
rect 9689 13277 9723 13311
rect 9965 13277 9999 13311
rect 4169 13209 4203 13243
rect 4629 13209 4663 13243
rect 7021 13209 7055 13243
rect 7205 13209 7239 13243
rect 7421 13209 7455 13243
rect 7665 13209 7699 13243
rect 7881 13209 7915 13243
rect 8493 13209 8527 13243
rect 1409 13141 1443 13175
rect 3157 13141 3191 13175
rect 3525 13141 3559 13175
rect 3801 13141 3835 13175
rect 3969 13141 4003 13175
rect 4905 13141 4939 13175
rect 8585 13141 8619 13175
rect 9873 13141 9907 13175
rect 13369 13141 13403 13175
rect 4353 12937 4387 12971
rect 6193 12937 6227 12971
rect 7205 12937 7239 12971
rect 7849 12937 7883 12971
rect 2881 12869 2915 12903
rect 6377 12869 6411 12903
rect 6593 12869 6627 12903
rect 8309 12869 8343 12903
rect 7021 12801 7055 12835
rect 7297 12801 7331 12835
rect 7665 12801 7699 12835
rect 7849 12801 7883 12835
rect 7941 12801 7975 12835
rect 10333 12801 10367 12835
rect 11989 12801 12023 12835
rect 2605 12733 2639 12767
rect 4445 12733 4479 12767
rect 4721 12733 4755 12767
rect 8033 12733 8067 12767
rect 6561 12597 6595 12631
rect 6745 12597 6779 12631
rect 6929 12597 6963 12631
rect 9781 12597 9815 12631
rect 10425 12597 10459 12631
rect 12081 12597 12115 12631
rect 4353 12393 4387 12427
rect 4813 12393 4847 12427
rect 6285 12393 6319 12427
rect 6469 12393 6503 12427
rect 8217 12393 8251 12427
rect 5549 12257 5583 12291
rect 9321 12257 9355 12291
rect 11161 12257 11195 12291
rect 4261 12189 4295 12223
rect 4445 12189 4479 12223
rect 5089 12189 5123 12223
rect 5181 12189 5215 12223
rect 5273 12189 5307 12223
rect 5457 12189 5491 12223
rect 5733 12189 5767 12223
rect 6009 12189 6043 12223
rect 8401 12189 8435 12223
rect 8677 12189 8711 12223
rect 5917 12121 5951 12155
rect 6101 12121 6135 12155
rect 6317 12121 6351 12155
rect 9597 12121 9631 12155
rect 11437 12121 11471 12155
rect 8585 12053 8619 12087
rect 11069 12053 11103 12087
rect 12909 12053 12943 12087
rect 10241 11849 10275 11883
rect 12173 11849 12207 11883
rect 3617 11781 3651 11815
rect 5977 11781 6011 11815
rect 6193 11781 6227 11815
rect 8953 11781 8987 11815
rect 3709 11713 3743 11747
rect 5733 11713 5767 11747
rect 6377 11713 6411 11747
rect 6561 11713 6595 11747
rect 7021 11713 7055 11747
rect 10885 11713 10919 11747
rect 11069 11713 11103 11747
rect 11529 11713 11563 11747
rect 11713 11713 11747 11747
rect 11805 11713 11839 11747
rect 11897 11713 11931 11747
rect 1685 11645 1719 11679
rect 1961 11645 1995 11679
rect 10977 11645 11011 11679
rect 3433 11509 3467 11543
rect 4261 11509 4295 11543
rect 5825 11509 5859 11543
rect 6009 11509 6043 11543
rect 6745 11509 6779 11543
rect 6929 11509 6963 11543
rect 2145 11305 2179 11339
rect 2605 11305 2639 11339
rect 3433 11305 3467 11339
rect 4721 11305 4755 11339
rect 6929 11305 6963 11339
rect 9689 11305 9723 11339
rect 10149 11305 10183 11339
rect 11805 11305 11839 11339
rect 12357 11305 12391 11339
rect 2421 11237 2455 11271
rect 5089 11237 5123 11271
rect 11069 11237 11103 11271
rect 5457 11169 5491 11203
rect 11345 11169 11379 11203
rect 11437 11169 11471 11203
rect 11620 11169 11654 11203
rect 2329 11101 2363 11135
rect 3249 11101 3283 11135
rect 3525 11101 3559 11135
rect 4637 11101 4671 11135
rect 4905 11101 4939 11135
rect 5181 11101 5215 11135
rect 10425 11101 10459 11135
rect 10517 11101 10551 11135
rect 10609 11101 10643 11135
rect 10793 11101 10827 11135
rect 10885 11101 10919 11135
rect 11539 11101 11573 11135
rect 11897 11101 11931 11135
rect 12265 11101 12299 11135
rect 12449 11101 12483 11135
rect 12541 11101 12575 11135
rect 2589 11033 2623 11067
rect 2789 11033 2823 11067
rect 3065 11033 3099 11067
rect 4077 11033 4111 11067
rect 9045 11033 9079 11067
rect 9873 11033 9907 11067
rect 11989 11033 12023 11067
rect 12173 11033 12207 11067
rect 2881 10965 2915 10999
rect 9505 10965 9539 10999
rect 9673 10965 9707 10999
rect 11897 10965 11931 10999
rect 12633 10965 12667 10999
rect 1685 10761 1719 10795
rect 4261 10761 4295 10795
rect 5089 10761 5123 10795
rect 7021 10761 7055 10795
rect 7665 10761 7699 10795
rect 7757 10761 7791 10795
rect 8585 10761 8619 10795
rect 2053 10693 2087 10727
rect 3801 10693 3835 10727
rect 4017 10693 4051 10727
rect 5701 10693 5735 10727
rect 5917 10693 5951 10727
rect 6837 10693 6871 10727
rect 9137 10693 9171 10727
rect 1501 10625 1535 10659
rect 4445 10625 4479 10659
rect 4997 10625 5031 10659
rect 5273 10625 5307 10659
rect 5365 10625 5399 10659
rect 6561 10625 6595 10659
rect 7389 10625 7423 10659
rect 7573 10625 7607 10659
rect 7941 10625 7975 10659
rect 8033 10625 8067 10659
rect 10701 10625 10735 10659
rect 10885 10625 10919 10659
rect 10977 10625 11011 10659
rect 11069 10625 11103 10659
rect 11529 10625 11563 10659
rect 1777 10557 1811 10591
rect 4629 10557 4663 10591
rect 6377 10557 6411 10591
rect 8677 10557 8711 10591
rect 9505 10557 9539 10591
rect 9597 10557 9631 10591
rect 9689 10557 9723 10591
rect 9781 10557 9815 10591
rect 11345 10557 11379 10591
rect 11805 10557 11839 10591
rect 4169 10489 4203 10523
rect 6745 10489 6779 10523
rect 8401 10489 8435 10523
rect 9137 10489 9171 10523
rect 3525 10421 3559 10455
rect 3985 10421 4019 10455
rect 4905 10421 4939 10455
rect 5549 10421 5583 10455
rect 5733 10421 5767 10455
rect 7021 10421 7055 10455
rect 7205 10421 7239 10455
rect 8217 10421 8251 10455
rect 9321 10421 9355 10455
rect 13277 10421 13311 10455
rect 2329 10217 2363 10251
rect 2513 10217 2547 10251
rect 2789 10217 2823 10251
rect 6745 10217 6779 10251
rect 8217 10217 8251 10251
rect 11161 10217 11195 10251
rect 11437 10217 11471 10251
rect 3893 10149 3927 10183
rect 12725 10149 12759 10183
rect 3617 10081 3651 10115
rect 4905 10081 4939 10115
rect 7389 10081 7423 10115
rect 11989 10081 12023 10115
rect 2973 10013 3007 10047
rect 3341 10013 3375 10047
rect 3433 10013 3467 10047
rect 3801 10013 3835 10047
rect 3985 10013 4019 10047
rect 4169 10013 4203 10047
rect 4353 10013 4387 10047
rect 4445 10013 4479 10047
rect 4537 10013 4571 10047
rect 7481 10013 7515 10047
rect 7849 10013 7883 10047
rect 8125 10013 8159 10047
rect 8309 10013 8343 10047
rect 8493 10013 8527 10047
rect 8585 10013 8619 10047
rect 8953 10013 8987 10047
rect 9137 10013 9171 10047
rect 9413 10013 9447 10047
rect 9689 10013 9723 10047
rect 11621 10013 11655 10047
rect 11713 10013 11747 10047
rect 12081 10013 12115 10047
rect 12357 10013 12391 10047
rect 2697 9945 2731 9979
rect 3157 9945 3191 9979
rect 4813 9945 4847 9979
rect 5181 9945 5215 9979
rect 7573 9945 7607 9979
rect 9597 9945 9631 9979
rect 10977 9945 11011 9979
rect 11193 9945 11227 9979
rect 12541 9945 12575 9979
rect 2497 9877 2531 9911
rect 6653 9877 6687 9911
rect 8033 9877 8067 9911
rect 8769 9877 8803 9911
rect 9321 9877 9355 9911
rect 11345 9877 11379 9911
rect 11805 9877 11839 9911
rect 12173 9877 12207 9911
rect 12449 9877 12483 9911
rect 4721 9673 4755 9707
rect 9689 9673 9723 9707
rect 2881 9605 2915 9639
rect 4537 9605 4571 9639
rect 4813 9605 4847 9639
rect 8217 9605 8251 9639
rect 2973 9537 3007 9571
rect 3249 9537 3283 9571
rect 4353 9537 4387 9571
rect 4445 9537 4479 9571
rect 5089 9537 5123 9571
rect 7941 9537 7975 9571
rect 11529 9537 11563 9571
rect 4905 9469 4939 9503
rect 11805 9469 11839 9503
rect 13277 9469 13311 9503
rect 4169 9401 4203 9435
rect 3157 9333 3191 9367
rect 4813 9333 4847 9367
rect 5273 9333 5307 9367
rect 2789 9129 2823 9163
rect 4077 9129 4111 9163
rect 4261 9129 4295 9163
rect 8401 9129 8435 9163
rect 8585 9129 8619 9163
rect 11069 9129 11103 9163
rect 12173 9129 12207 9163
rect 8217 8993 8251 9027
rect 11437 8993 11471 9027
rect 11621 8993 11655 9027
rect 11713 8993 11747 9027
rect 11897 8993 11931 9027
rect 12633 8993 12667 9027
rect 13277 8993 13311 9027
rect 2421 8925 2455 8959
rect 5273 8925 5307 8959
rect 5365 8925 5399 8959
rect 5549 8925 5583 8959
rect 5641 8925 5675 8959
rect 6561 8925 6595 8959
rect 10425 8925 10459 8959
rect 10609 8925 10643 8959
rect 10701 8925 10735 8959
rect 10793 8925 10827 8959
rect 11805 8925 11839 8959
rect 12081 8925 12115 8959
rect 2973 8857 3007 8891
rect 3893 8857 3927 8891
rect 4109 8857 4143 8891
rect 8769 8857 8803 8891
rect 2237 8789 2271 8823
rect 2605 8789 2639 8823
rect 2773 8789 2807 8823
rect 5825 8789 5859 8823
rect 8569 8789 8603 8823
rect 3433 8585 3467 8619
rect 3525 8585 3559 8619
rect 7665 8585 7699 8619
rect 8309 8585 8343 8619
rect 1961 8517 1995 8551
rect 3709 8517 3743 8551
rect 7817 8517 7851 8551
rect 7987 8517 8021 8551
rect 8861 8517 8895 8551
rect 1685 8449 1719 8483
rect 3893 8449 3927 8483
rect 6745 8449 6779 8483
rect 6837 8449 6871 8483
rect 7113 8449 7147 8483
rect 7297 8449 7331 8483
rect 8125 8449 8159 8483
rect 8217 8449 8251 8483
rect 8585 8449 8619 8483
rect 8677 8449 8711 8483
rect 10517 8449 10551 8483
rect 10701 8449 10735 8483
rect 6653 8381 6687 8415
rect 7021 8381 7055 8415
rect 8493 8381 8527 8415
rect 8401 8313 8435 8347
rect 7297 8245 7331 8279
rect 7889 8245 7923 8279
rect 8861 8245 8895 8279
rect 10609 8245 10643 8279
rect 2789 8041 2823 8075
rect 4721 8041 4755 8075
rect 4353 7973 4387 8007
rect 4905 7973 4939 8007
rect 4997 7973 5031 8007
rect 7941 7973 7975 8007
rect 10057 7973 10091 8007
rect 10517 7905 10551 7939
rect 10793 7905 10827 7939
rect 10977 7905 11011 7939
rect 2881 7837 2915 7871
rect 5181 7837 5215 7871
rect 5273 7837 5307 7871
rect 5457 7837 5491 7871
rect 8125 7837 8159 7871
rect 8585 7837 8619 7871
rect 8769 7837 8803 7871
rect 9689 7837 9723 7871
rect 9965 7837 9999 7871
rect 10149 7837 10183 7871
rect 10241 7837 10275 7871
rect 10425 7837 10459 7871
rect 10701 7837 10735 7871
rect 10885 7837 10919 7871
rect 11345 7837 11379 7871
rect 11437 7837 11471 7871
rect 11713 7837 11747 7871
rect 8217 7769 8251 7803
rect 8677 7769 8711 7803
rect 9597 7769 9631 7803
rect 11621 7769 11655 7803
rect 4721 7701 4755 7735
rect 5641 7701 5675 7735
rect 8309 7701 8343 7735
rect 8493 7701 8527 7735
rect 9781 7701 9815 7735
rect 11253 7701 11287 7735
rect 11713 7701 11747 7735
rect 4353 7497 4387 7531
rect 6469 7497 6503 7531
rect 6929 7497 6963 7531
rect 11621 7497 11655 7531
rect 11989 7497 12023 7531
rect 12281 7497 12315 7531
rect 12449 7497 12483 7531
rect 2973 7429 3007 7463
rect 4077 7429 4111 7463
rect 5917 7429 5951 7463
rect 8677 7429 8711 7463
rect 9781 7429 9815 7463
rect 12081 7429 12115 7463
rect 3157 7361 3191 7395
rect 3525 7361 3559 7395
rect 3985 7361 4019 7395
rect 4169 7361 4203 7395
rect 6561 7361 6595 7395
rect 6837 7361 6871 7395
rect 8033 7361 8067 7395
rect 8861 7361 8895 7395
rect 8953 7361 8987 7395
rect 9137 7361 9171 7395
rect 11529 7361 11563 7395
rect 11805 7361 11839 7395
rect 12725 7361 12759 7395
rect 13001 7361 13035 7395
rect 13093 7361 13127 7395
rect 3709 7293 3743 7327
rect 6193 7293 6227 7327
rect 8309 7293 8343 7327
rect 9045 7293 9079 7327
rect 9505 7293 9539 7327
rect 11253 7293 11287 7327
rect 3801 7225 3835 7259
rect 2789 7157 2823 7191
rect 3341 7157 3375 7191
rect 4445 7157 4479 7191
rect 12265 7157 12299 7191
rect 12541 7157 12575 7191
rect 12909 7157 12943 7191
rect 13185 7157 13219 7191
rect 2329 6953 2363 6987
rect 2789 6953 2823 6987
rect 7284 6953 7318 6987
rect 10425 6953 10459 6987
rect 11792 6953 11826 6987
rect 2145 6885 2179 6919
rect 2605 6885 2639 6919
rect 3249 6817 3283 6851
rect 4077 6817 4111 6851
rect 6653 6817 6687 6851
rect 7021 6817 7055 6851
rect 11529 6817 11563 6851
rect 13277 6817 13311 6851
rect 1869 6749 1903 6783
rect 2053 6749 2087 6783
rect 3157 6749 3191 6783
rect 3341 6749 3375 6783
rect 3433 6749 3467 6783
rect 3801 6749 3835 6783
rect 3985 6749 4019 6783
rect 6101 6749 6135 6783
rect 6929 6749 6963 6783
rect 9229 6749 9263 6783
rect 10057 6749 10091 6783
rect 10149 6749 10183 6783
rect 10793 6749 10827 6783
rect 10885 6749 10919 6783
rect 11253 6749 11287 6783
rect 2513 6681 2547 6715
rect 2973 6681 3007 6715
rect 4353 6681 4387 6715
rect 6009 6681 6043 6715
rect 9781 6681 9815 6715
rect 10517 6681 10551 6715
rect 11161 6681 11195 6715
rect 2053 6613 2087 6647
rect 2303 6613 2337 6647
rect 2773 6613 2807 6647
rect 3617 6613 3651 6647
rect 3985 6613 4019 6647
rect 5825 6613 5859 6647
rect 8769 6613 8803 6647
rect 9873 6613 9907 6647
rect 10609 6613 10643 6647
rect 11069 6613 11103 6647
rect 4445 6409 4479 6443
rect 5089 6409 5123 6443
rect 6653 6409 6687 6443
rect 8217 6409 8251 6443
rect 9505 6409 9539 6443
rect 9781 6409 9815 6443
rect 10625 6409 10659 6443
rect 11253 6409 11287 6443
rect 13277 6409 13311 6443
rect 10425 6341 10459 6375
rect 1501 6273 1535 6307
rect 1777 6273 1811 6307
rect 3801 6273 3835 6307
rect 3985 6273 4019 6307
rect 4077 6273 4111 6307
rect 4169 6273 4203 6307
rect 4629 6273 4663 6307
rect 4813 6273 4847 6307
rect 6469 6273 6503 6307
rect 8033 6273 8067 6307
rect 8125 6273 8159 6307
rect 8677 6273 8711 6307
rect 9137 6273 9171 6307
rect 9229 6273 9263 6307
rect 9597 6273 9631 6307
rect 9689 6259 9723 6293
rect 9789 6271 9823 6305
rect 9965 6273 9999 6307
rect 10057 6273 10091 6307
rect 10885 6273 10919 6307
rect 11069 6273 11103 6307
rect 11345 6273 11379 6307
rect 2053 6205 2087 6239
rect 4721 6205 4755 6239
rect 4905 6205 4939 6239
rect 7849 6205 7883 6239
rect 8769 6205 8803 6239
rect 11529 6205 11563 6239
rect 11805 6205 11839 6239
rect 1685 6137 1719 6171
rect 10977 6137 11011 6171
rect 3525 6069 3559 6103
rect 8493 6069 8527 6103
rect 9045 6069 9079 6103
rect 10149 6069 10183 6103
rect 10609 6069 10643 6103
rect 10793 6069 10827 6103
rect 3801 5865 3835 5899
rect 5273 5865 5307 5899
rect 10425 5865 10459 5899
rect 11345 5865 11379 5899
rect 3249 5797 3283 5831
rect 1501 5729 1535 5763
rect 3525 5729 3559 5763
rect 3617 5661 3651 5695
rect 3985 5661 4019 5695
rect 6561 5661 6595 5695
rect 9137 5661 9171 5695
rect 11161 5661 11195 5695
rect 1777 5593 1811 5627
rect 4169 5593 4203 5627
rect 2145 5321 2179 5355
rect 2973 5321 3007 5355
rect 3249 5253 3283 5287
rect 4905 5253 4939 5287
rect 2329 5185 2363 5219
rect 3065 5185 3099 5219
rect 3341 5185 3375 5219
rect 5549 5117 5583 5151
rect 5917 5049 5951 5083
rect 6009 4981 6043 5015
rect 4813 4777 4847 4811
rect 7205 4709 7239 4743
rect 5457 4641 5491 4675
rect 9413 4641 9447 4675
rect 9597 4641 9631 4675
rect 10333 4641 10367 4675
rect 4353 4573 4387 4607
rect 7481 4573 7515 4607
rect 8401 4573 8435 4607
rect 8953 4573 8987 4607
rect 9505 4573 9539 4607
rect 9689 4573 9723 4607
rect 10057 4573 10091 4607
rect 12633 4573 12667 4607
rect 13093 4573 13127 4607
rect 4997 4505 5031 4539
rect 5733 4505 5767 4539
rect 7389 4505 7423 4539
rect 8585 4505 8619 4539
rect 10609 4505 10643 4539
rect 4169 4437 4203 4471
rect 4629 4437 4663 4471
rect 4797 4437 4831 4471
rect 8769 4437 8803 4471
rect 9137 4437 9171 4471
rect 9229 4437 9263 4471
rect 10241 4437 10275 4471
rect 12081 4437 12115 4471
rect 12541 4437 12575 4471
rect 13277 4437 13311 4471
rect 4261 4233 4295 4267
rect 5825 4233 5859 4267
rect 10793 4233 10827 4267
rect 10977 4233 11011 4267
rect 4077 4165 4111 4199
rect 5457 4165 5491 4199
rect 5641 4165 5675 4199
rect 6529 4165 6563 4199
rect 6745 4165 6779 4199
rect 6929 4165 6963 4199
rect 10885 4165 10919 4199
rect 4629 4097 4663 4131
rect 4813 4097 4847 4131
rect 5273 4097 5307 4131
rect 5365 4097 5399 4131
rect 6009 4097 6043 4131
rect 6837 4097 6871 4131
rect 7021 4097 7055 4131
rect 9781 4097 9815 4131
rect 10057 4097 10091 4131
rect 10517 4097 10551 4131
rect 10609 4097 10643 4131
rect 11897 4097 11931 4131
rect 12265 4097 12299 4131
rect 13001 4097 13035 4131
rect 13093 4097 13127 4131
rect 4353 4029 4387 4063
rect 4537 4029 4571 4063
rect 4721 4029 4755 4063
rect 9505 4029 9539 4063
rect 10149 4029 10183 4063
rect 11805 4029 11839 4063
rect 12817 4029 12851 4063
rect 3709 3961 3743 3995
rect 4077 3893 4111 3927
rect 5089 3893 5123 3927
rect 6377 3893 6411 3927
rect 6561 3893 6595 3927
rect 8033 3893 8067 3927
rect 9873 3893 9907 3927
rect 10057 3893 10091 3927
rect 11161 3893 11195 3927
rect 11529 3893 11563 3927
rect 5549 3689 5583 3723
rect 7665 3689 7699 3723
rect 8677 3689 8711 3723
rect 9210 3689 9244 3723
rect 10701 3689 10735 3723
rect 12541 3689 12575 3723
rect 1409 3621 1443 3655
rect 3801 3553 3835 3587
rect 5917 3553 5951 3587
rect 8493 3553 8527 3587
rect 8953 3553 8987 3587
rect 10793 3553 10827 3587
rect 11069 3553 11103 3587
rect 3157 3485 3191 3519
rect 3433 3485 3467 3519
rect 5641 3485 5675 3519
rect 7941 3485 7975 3519
rect 8401 3485 8435 3519
rect 13369 3485 13403 3519
rect 4077 3417 4111 3451
rect 6193 3417 6227 3451
rect 8033 3417 8067 3451
rect 3341 3349 3375 3383
rect 3525 3349 3559 3383
rect 5825 3349 5859 3383
rect 4997 3145 5031 3179
rect 5365 3145 5399 3179
rect 5825 3145 5859 3179
rect 6377 3145 6411 3179
rect 7021 3145 7055 3179
rect 8309 3145 8343 3179
rect 8693 3145 8727 3179
rect 8861 3145 8895 3179
rect 9321 3145 9355 3179
rect 9505 3145 9539 3179
rect 5549 3077 5583 3111
rect 6745 3077 6779 3111
rect 8493 3077 8527 3111
rect 3157 3009 3191 3043
rect 5181 3009 5215 3043
rect 5457 3009 5491 3043
rect 5733 3009 5767 3043
rect 5825 3009 5859 3043
rect 6561 3009 6595 3043
rect 6929 3009 6963 3043
rect 8217 3009 8251 3043
rect 9597 3009 9631 3043
rect 1409 2941 1443 2975
rect 3433 2941 3467 2975
rect 4905 2941 4939 2975
rect 8953 2941 8987 2975
rect 10241 2941 10275 2975
rect 13369 2941 13403 2975
rect 8677 2805 8711 2839
rect 9321 2805 9355 2839
rect 4169 2601 4203 2635
rect 7389 2601 7423 2635
rect 4077 2397 4111 2431
rect 7205 2397 7239 2431
rect 9413 2397 9447 2431
rect 10057 2397 10091 2431
rect 10701 2397 10735 2431
rect 9229 2261 9263 2295
rect 9873 2261 9907 2295
rect 10517 2261 10551 2295
<< metal1 >>
rect 1104 14714 13708 14736
rect 1104 14662 2525 14714
rect 2577 14662 2589 14714
rect 2641 14662 2653 14714
rect 2705 14662 2717 14714
rect 2769 14662 2781 14714
rect 2833 14662 5676 14714
rect 5728 14662 5740 14714
rect 5792 14662 5804 14714
rect 5856 14662 5868 14714
rect 5920 14662 5932 14714
rect 5984 14662 8827 14714
rect 8879 14662 8891 14714
rect 8943 14662 8955 14714
rect 9007 14662 9019 14714
rect 9071 14662 9083 14714
rect 9135 14662 11978 14714
rect 12030 14662 12042 14714
rect 12094 14662 12106 14714
rect 12158 14662 12170 14714
rect 12222 14662 12234 14714
rect 12286 14662 13708 14714
rect 1104 14640 13708 14662
rect 1104 14170 13708 14192
rect 1104 14118 3185 14170
rect 3237 14118 3249 14170
rect 3301 14118 3313 14170
rect 3365 14118 3377 14170
rect 3429 14118 3441 14170
rect 3493 14118 6336 14170
rect 6388 14118 6400 14170
rect 6452 14118 6464 14170
rect 6516 14118 6528 14170
rect 6580 14118 6592 14170
rect 6644 14118 9487 14170
rect 9539 14118 9551 14170
rect 9603 14118 9615 14170
rect 9667 14118 9679 14170
rect 9731 14118 9743 14170
rect 9795 14118 12638 14170
rect 12690 14118 12702 14170
rect 12754 14118 12766 14170
rect 12818 14118 12830 14170
rect 12882 14118 12894 14170
rect 12946 14118 13708 14170
rect 1104 14096 13708 14118
rect 9582 13988 9588 14000
rect 9062 13960 9588 13988
rect 9582 13948 9588 13960
rect 9640 13948 9646 14000
rect 5721 13923 5779 13929
rect 5721 13889 5733 13923
rect 5767 13920 5779 13923
rect 6454 13920 6460 13932
rect 5767 13892 6460 13920
rect 5767 13889 5779 13892
rect 5721 13883 5779 13889
rect 6454 13880 6460 13892
rect 6512 13880 6518 13932
rect 6549 13923 6607 13929
rect 6549 13889 6561 13923
rect 6595 13920 6607 13923
rect 6730 13920 6736 13932
rect 6595 13892 6736 13920
rect 6595 13889 6607 13892
rect 6549 13883 6607 13889
rect 6730 13880 6736 13892
rect 6788 13880 6794 13932
rect 1394 13812 1400 13864
rect 1452 13812 1458 13864
rect 5810 13812 5816 13864
rect 5868 13812 5874 13864
rect 5905 13855 5963 13861
rect 5905 13821 5917 13855
rect 5951 13821 5963 13855
rect 5905 13815 5963 13821
rect 5997 13855 6055 13861
rect 5997 13821 6009 13855
rect 6043 13821 6055 13855
rect 5997 13815 6055 13821
rect 5534 13744 5540 13796
rect 5592 13784 5598 13796
rect 5920 13784 5948 13815
rect 5592 13756 5948 13784
rect 5592 13744 5598 13756
rect 4614 13676 4620 13728
rect 4672 13716 4678 13728
rect 5442 13716 5448 13728
rect 4672 13688 5448 13716
rect 4672 13676 4678 13688
rect 5442 13676 5448 13688
rect 5500 13716 5506 13728
rect 6012 13716 6040 13815
rect 9490 13812 9496 13864
rect 9548 13812 9554 13864
rect 9769 13855 9827 13861
rect 9769 13821 9781 13855
rect 9815 13852 9827 13855
rect 10226 13852 10232 13864
rect 9815 13824 10232 13852
rect 9815 13821 9827 13824
rect 9769 13815 9827 13821
rect 10226 13812 10232 13824
rect 10284 13812 10290 13864
rect 13354 13812 13360 13864
rect 13412 13812 13418 13864
rect 5500 13688 6040 13716
rect 5500 13676 5506 13688
rect 6178 13676 6184 13728
rect 6236 13676 6242 13728
rect 6362 13676 6368 13728
rect 6420 13676 6426 13728
rect 7926 13676 7932 13728
rect 7984 13716 7990 13728
rect 8021 13719 8079 13725
rect 8021 13716 8033 13719
rect 7984 13688 8033 13716
rect 7984 13676 7990 13688
rect 8021 13685 8033 13688
rect 8067 13685 8079 13719
rect 8021 13679 8079 13685
rect 1104 13626 13708 13648
rect 1104 13574 2525 13626
rect 2577 13574 2589 13626
rect 2641 13574 2653 13626
rect 2705 13574 2717 13626
rect 2769 13574 2781 13626
rect 2833 13574 5676 13626
rect 5728 13574 5740 13626
rect 5792 13574 5804 13626
rect 5856 13574 5868 13626
rect 5920 13574 5932 13626
rect 5984 13574 8827 13626
rect 8879 13574 8891 13626
rect 8943 13574 8955 13626
rect 9007 13574 9019 13626
rect 9071 13574 9083 13626
rect 9135 13574 11978 13626
rect 12030 13574 12042 13626
rect 12094 13574 12106 13626
rect 12158 13574 12170 13626
rect 12222 13574 12234 13626
rect 12286 13574 13708 13626
rect 1104 13552 13708 13574
rect 3973 13515 4031 13521
rect 3973 13481 3985 13515
rect 4019 13512 4031 13515
rect 4249 13515 4307 13521
rect 4249 13512 4261 13515
rect 4019 13484 4261 13512
rect 4019 13481 4031 13484
rect 3973 13475 4031 13481
rect 4249 13481 4261 13484
rect 4295 13481 4307 13515
rect 4249 13475 4307 13481
rect 4798 13472 4804 13524
rect 4856 13512 4862 13524
rect 5994 13512 6000 13524
rect 4856 13484 6000 13512
rect 4856 13472 4862 13484
rect 5994 13472 6000 13484
rect 6052 13472 6058 13524
rect 6454 13472 6460 13524
rect 6512 13512 6518 13524
rect 6822 13512 6828 13524
rect 6512 13484 6828 13512
rect 6512 13472 6518 13484
rect 6822 13472 6828 13484
rect 6880 13472 6886 13524
rect 7377 13515 7435 13521
rect 7377 13481 7389 13515
rect 7423 13512 7435 13515
rect 7423 13484 7788 13512
rect 7423 13481 7435 13484
rect 7377 13475 7435 13481
rect 7561 13447 7619 13453
rect 7561 13413 7573 13447
rect 7607 13413 7619 13447
rect 7760 13444 7788 13484
rect 7834 13472 7840 13524
rect 7892 13472 7898 13524
rect 9033 13515 9091 13521
rect 9033 13512 9045 13515
rect 7944 13484 9045 13512
rect 7944 13444 7972 13484
rect 9033 13481 9045 13484
rect 9079 13481 9091 13515
rect 9033 13475 9091 13481
rect 9401 13515 9459 13521
rect 9401 13481 9413 13515
rect 9447 13512 9459 13515
rect 9490 13512 9496 13524
rect 9447 13484 9496 13512
rect 9447 13481 9459 13484
rect 9401 13475 9459 13481
rect 9490 13472 9496 13484
rect 9548 13472 9554 13524
rect 9582 13472 9588 13524
rect 9640 13472 9646 13524
rect 7760 13416 7972 13444
rect 8021 13447 8079 13453
rect 7561 13407 7619 13413
rect 8021 13413 8033 13447
rect 8067 13444 8079 13447
rect 8067 13416 9260 13444
rect 8067 13413 8079 13416
rect 8021 13407 8079 13413
rect 4154 13336 4160 13388
rect 4212 13376 4218 13388
rect 5077 13379 5135 13385
rect 5077 13376 5089 13379
rect 4212 13348 5089 13376
rect 4212 13336 4218 13348
rect 5077 13345 5089 13348
rect 5123 13345 5135 13379
rect 5077 13339 5135 13345
rect 5353 13379 5411 13385
rect 5353 13345 5365 13379
rect 5399 13376 5411 13379
rect 6362 13376 6368 13388
rect 5399 13348 6368 13376
rect 5399 13345 5411 13348
rect 5353 13339 5411 13345
rect 6362 13336 6368 13348
rect 6420 13336 6426 13388
rect 7576 13376 7604 13407
rect 7576 13348 8800 13376
rect 3329 13311 3387 13317
rect 3329 13277 3341 13311
rect 3375 13277 3387 13311
rect 3329 13271 3387 13277
rect 3421 13311 3479 13317
rect 3421 13277 3433 13311
rect 3467 13308 3479 13311
rect 3694 13308 3700 13320
rect 3467 13280 3700 13308
rect 3467 13277 3479 13280
rect 3421 13271 3479 13277
rect 3344 13240 3372 13271
rect 3694 13268 3700 13280
rect 3752 13268 3758 13320
rect 4433 13311 4491 13317
rect 4433 13277 4445 13311
rect 4479 13308 4491 13311
rect 4798 13308 4804 13320
rect 4479 13280 4804 13308
rect 4479 13277 4491 13280
rect 4433 13271 4491 13277
rect 4798 13268 4804 13280
rect 4856 13268 4862 13320
rect 4985 13311 5043 13317
rect 4985 13277 4997 13311
rect 5031 13277 5043 13311
rect 4985 13271 5043 13277
rect 4157 13243 4215 13249
rect 3344 13212 3832 13240
rect 842 13132 848 13184
rect 900 13172 906 13184
rect 1397 13175 1455 13181
rect 1397 13172 1409 13175
rect 900 13144 1409 13172
rect 900 13132 906 13144
rect 1397 13141 1409 13144
rect 1443 13141 1455 13175
rect 1397 13135 1455 13141
rect 2866 13132 2872 13184
rect 2924 13172 2930 13184
rect 3145 13175 3203 13181
rect 3145 13172 3157 13175
rect 2924 13144 3157 13172
rect 2924 13132 2930 13144
rect 3145 13141 3157 13144
rect 3191 13141 3203 13175
rect 3145 13135 3203 13141
rect 3510 13132 3516 13184
rect 3568 13132 3574 13184
rect 3804 13181 3832 13212
rect 4157 13209 4169 13243
rect 4203 13240 4215 13243
rect 4522 13240 4528 13252
rect 4203 13212 4528 13240
rect 4203 13209 4215 13212
rect 4157 13203 4215 13209
rect 4522 13200 4528 13212
rect 4580 13200 4586 13252
rect 4614 13200 4620 13252
rect 4672 13200 4678 13252
rect 5000 13240 5028 13271
rect 7098 13268 7104 13320
rect 7156 13268 7162 13320
rect 8113 13311 8171 13317
rect 8113 13308 8125 13311
rect 7576 13280 8125 13308
rect 7009 13243 7067 13249
rect 7009 13240 7021 13243
rect 5000 13212 5580 13240
rect 6578 13212 7021 13240
rect 5552 13184 5580 13212
rect 7009 13209 7021 13212
rect 7055 13209 7067 13243
rect 7009 13203 7067 13209
rect 7190 13200 7196 13252
rect 7248 13200 7254 13252
rect 7409 13243 7467 13249
rect 7409 13209 7421 13243
rect 7455 13240 7467 13243
rect 7576 13240 7604 13280
rect 8113 13277 8125 13280
rect 8159 13277 8171 13311
rect 8113 13271 8171 13277
rect 8297 13311 8355 13317
rect 8297 13277 8309 13311
rect 8343 13308 8355 13311
rect 8386 13308 8392 13320
rect 8343 13280 8392 13308
rect 8343 13277 8355 13280
rect 8297 13271 8355 13277
rect 8386 13268 8392 13280
rect 8444 13308 8450 13320
rect 8772 13317 8800 13348
rect 8757 13311 8815 13317
rect 8444 13280 8708 13308
rect 8444 13268 8450 13280
rect 7455 13212 7604 13240
rect 7653 13243 7711 13249
rect 7455 13209 7467 13212
rect 7409 13203 7467 13209
rect 7653 13209 7665 13243
rect 7699 13209 7711 13243
rect 7653 13203 7711 13209
rect 7869 13243 7927 13249
rect 7869 13209 7881 13243
rect 7915 13240 7927 13243
rect 8202 13240 8208 13252
rect 7915 13212 8208 13240
rect 7915 13209 7927 13212
rect 7869 13203 7927 13209
rect 3789 13175 3847 13181
rect 3789 13141 3801 13175
rect 3835 13141 3847 13175
rect 3789 13135 3847 13141
rect 3957 13175 4015 13181
rect 3957 13141 3969 13175
rect 4003 13172 4015 13175
rect 4338 13172 4344 13184
rect 4003 13144 4344 13172
rect 4003 13141 4015 13144
rect 3957 13135 4015 13141
rect 4338 13132 4344 13144
rect 4396 13132 4402 13184
rect 4893 13175 4951 13181
rect 4893 13141 4905 13175
rect 4939 13172 4951 13175
rect 5074 13172 5080 13184
rect 4939 13144 5080 13172
rect 4939 13141 4951 13144
rect 4893 13135 4951 13141
rect 5074 13132 5080 13144
rect 5132 13132 5138 13184
rect 5534 13132 5540 13184
rect 5592 13132 5598 13184
rect 7208 13172 7236 13200
rect 7668 13172 7696 13203
rect 8202 13200 8208 13212
rect 8260 13200 8266 13252
rect 8478 13200 8484 13252
rect 8536 13200 8542 13252
rect 8680 13240 8708 13280
rect 8757 13277 8769 13311
rect 8803 13277 8815 13311
rect 8757 13271 8815 13277
rect 8941 13311 8999 13317
rect 8941 13277 8953 13311
rect 8987 13277 8999 13311
rect 8941 13271 8999 13277
rect 8956 13240 8984 13271
rect 9122 13268 9128 13320
rect 9180 13268 9186 13320
rect 9232 13317 9260 13416
rect 9217 13311 9275 13317
rect 9217 13277 9229 13311
rect 9263 13277 9275 13311
rect 9217 13271 9275 13277
rect 9677 13311 9735 13317
rect 9677 13277 9689 13311
rect 9723 13308 9735 13311
rect 9953 13311 10011 13317
rect 9953 13308 9965 13311
rect 9723 13280 9965 13308
rect 9723 13277 9735 13280
rect 9677 13271 9735 13277
rect 9953 13277 9965 13280
rect 9999 13308 10011 13311
rect 10410 13308 10416 13320
rect 9999 13280 10416 13308
rect 9999 13277 10011 13280
rect 9953 13271 10011 13277
rect 10410 13268 10416 13280
rect 10468 13268 10474 13320
rect 9398 13240 9404 13252
rect 8680 13212 9404 13240
rect 9398 13200 9404 13212
rect 9456 13200 9462 13252
rect 7208 13144 7696 13172
rect 7742 13132 7748 13184
rect 7800 13172 7806 13184
rect 8496 13172 8524 13200
rect 7800 13144 8524 13172
rect 7800 13132 7806 13144
rect 8570 13132 8576 13184
rect 8628 13132 8634 13184
rect 9858 13132 9864 13184
rect 9916 13132 9922 13184
rect 13354 13132 13360 13184
rect 13412 13132 13418 13184
rect 1104 13082 13708 13104
rect 1104 13030 3185 13082
rect 3237 13030 3249 13082
rect 3301 13030 3313 13082
rect 3365 13030 3377 13082
rect 3429 13030 3441 13082
rect 3493 13030 6336 13082
rect 6388 13030 6400 13082
rect 6452 13030 6464 13082
rect 6516 13030 6528 13082
rect 6580 13030 6592 13082
rect 6644 13030 9487 13082
rect 9539 13030 9551 13082
rect 9603 13030 9615 13082
rect 9667 13030 9679 13082
rect 9731 13030 9743 13082
rect 9795 13030 12638 13082
rect 12690 13030 12702 13082
rect 12754 13030 12766 13082
rect 12818 13030 12830 13082
rect 12882 13030 12894 13082
rect 12946 13030 13708 13082
rect 1104 13008 13708 13030
rect 4341 12971 4399 12977
rect 4341 12937 4353 12971
rect 4387 12968 4399 12971
rect 4798 12968 4804 12980
rect 4387 12940 4804 12968
rect 4387 12937 4399 12940
rect 4341 12931 4399 12937
rect 4798 12928 4804 12940
rect 4856 12928 4862 12980
rect 5534 12928 5540 12980
rect 5592 12968 5598 12980
rect 6086 12968 6092 12980
rect 5592 12940 6092 12968
rect 5592 12928 5598 12940
rect 6086 12928 6092 12940
rect 6144 12968 6150 12980
rect 6181 12971 6239 12977
rect 6181 12968 6193 12971
rect 6144 12940 6193 12968
rect 6144 12928 6150 12940
rect 6181 12937 6193 12940
rect 6227 12937 6239 12971
rect 7193 12971 7251 12977
rect 7193 12968 7205 12971
rect 6181 12931 6239 12937
rect 6288 12940 7205 12968
rect 2866 12860 2872 12912
rect 2924 12860 2930 12912
rect 3510 12860 3516 12912
rect 3568 12860 3574 12912
rect 6288 12900 6316 12940
rect 7193 12937 7205 12940
rect 7239 12937 7251 12971
rect 7193 12931 7251 12937
rect 7834 12928 7840 12980
rect 7892 12928 7898 12980
rect 8386 12968 8392 12980
rect 8220 12940 8392 12968
rect 5934 12872 6316 12900
rect 6365 12903 6423 12909
rect 6365 12869 6377 12903
rect 6411 12869 6423 12903
rect 6365 12863 6423 12869
rect 6581 12903 6639 12909
rect 6581 12869 6593 12903
rect 6627 12900 6639 12903
rect 6822 12900 6828 12912
rect 6627 12872 6828 12900
rect 6627 12869 6639 12872
rect 6581 12863 6639 12869
rect 5994 12792 6000 12844
rect 6052 12832 6058 12844
rect 6380 12832 6408 12863
rect 6822 12860 6828 12872
rect 6880 12860 6886 12912
rect 8220 12900 8248 12940
rect 8386 12928 8392 12940
rect 8444 12928 8450 12980
rect 8478 12928 8484 12980
rect 8536 12968 8542 12980
rect 9122 12968 9128 12980
rect 8536 12940 9128 12968
rect 8536 12928 8542 12940
rect 9122 12928 9128 12940
rect 9180 12928 9186 12980
rect 7852 12872 8248 12900
rect 8297 12903 8355 12909
rect 6052 12804 6408 12832
rect 7009 12835 7067 12841
rect 6052 12792 6058 12804
rect 7009 12801 7021 12835
rect 7055 12801 7067 12835
rect 7009 12795 7067 12801
rect 1670 12724 1676 12776
rect 1728 12764 1734 12776
rect 2593 12767 2651 12773
rect 2593 12764 2605 12767
rect 1728 12736 2605 12764
rect 1728 12724 1734 12736
rect 2593 12733 2605 12736
rect 2639 12733 2651 12767
rect 2593 12727 2651 12733
rect 4154 12724 4160 12776
rect 4212 12764 4218 12776
rect 4433 12767 4491 12773
rect 4433 12764 4445 12767
rect 4212 12736 4445 12764
rect 4212 12724 4218 12736
rect 4433 12733 4445 12736
rect 4479 12733 4491 12767
rect 4433 12727 4491 12733
rect 4706 12724 4712 12776
rect 4764 12724 4770 12776
rect 7024 12764 7052 12795
rect 7098 12792 7104 12844
rect 7156 12832 7162 12844
rect 7285 12835 7343 12841
rect 7285 12832 7297 12835
rect 7156 12804 7297 12832
rect 7156 12792 7162 12804
rect 7285 12801 7297 12804
rect 7331 12801 7343 12835
rect 7285 12795 7343 12801
rect 7653 12835 7711 12841
rect 7653 12801 7665 12835
rect 7699 12832 7711 12835
rect 7742 12832 7748 12844
rect 7699 12804 7748 12832
rect 7699 12801 7711 12804
rect 7653 12795 7711 12801
rect 7668 12764 7696 12795
rect 7742 12792 7748 12804
rect 7800 12792 7806 12844
rect 7852 12841 7880 12872
rect 8297 12869 8309 12903
rect 8343 12900 8355 12903
rect 8570 12900 8576 12912
rect 8343 12872 8576 12900
rect 8343 12869 8355 12872
rect 8297 12863 8355 12869
rect 8570 12860 8576 12872
rect 8628 12860 8634 12912
rect 9858 12900 9864 12912
rect 9522 12872 9864 12900
rect 9858 12860 9864 12872
rect 9916 12860 9922 12912
rect 7837 12835 7895 12841
rect 7837 12801 7849 12835
rect 7883 12801 7895 12835
rect 7837 12795 7895 12801
rect 7926 12792 7932 12844
rect 7984 12792 7990 12844
rect 10321 12835 10379 12841
rect 10321 12801 10333 12835
rect 10367 12832 10379 12835
rect 10410 12832 10416 12844
rect 10367 12804 10416 12832
rect 10367 12801 10379 12804
rect 10321 12795 10379 12801
rect 10410 12792 10416 12804
rect 10468 12832 10474 12844
rect 11977 12835 12035 12841
rect 11977 12832 11989 12835
rect 10468 12804 11989 12832
rect 10468 12792 10474 12804
rect 11977 12801 11989 12804
rect 12023 12801 12035 12835
rect 11977 12795 12035 12801
rect 7024 12736 7696 12764
rect 8021 12767 8079 12773
rect 8021 12733 8033 12767
rect 8067 12733 8079 12767
rect 8021 12727 8079 12733
rect 7926 12656 7932 12708
rect 7984 12696 7990 12708
rect 8036 12696 8064 12727
rect 7984 12668 8064 12696
rect 7984 12656 7990 12668
rect 6086 12588 6092 12640
rect 6144 12628 6150 12640
rect 6549 12631 6607 12637
rect 6549 12628 6561 12631
rect 6144 12600 6561 12628
rect 6144 12588 6150 12600
rect 6549 12597 6561 12600
rect 6595 12597 6607 12631
rect 6549 12591 6607 12597
rect 6733 12631 6791 12637
rect 6733 12597 6745 12631
rect 6779 12628 6791 12631
rect 6822 12628 6828 12640
rect 6779 12600 6828 12628
rect 6779 12597 6791 12600
rect 6733 12591 6791 12597
rect 6822 12588 6828 12600
rect 6880 12588 6886 12640
rect 6914 12588 6920 12640
rect 6972 12588 6978 12640
rect 8018 12588 8024 12640
rect 8076 12628 8082 12640
rect 8386 12628 8392 12640
rect 8076 12600 8392 12628
rect 8076 12588 8082 12600
rect 8386 12588 8392 12600
rect 8444 12588 8450 12640
rect 9398 12588 9404 12640
rect 9456 12628 9462 12640
rect 9769 12631 9827 12637
rect 9769 12628 9781 12631
rect 9456 12600 9781 12628
rect 9456 12588 9462 12600
rect 9769 12597 9781 12600
rect 9815 12597 9827 12631
rect 9769 12591 9827 12597
rect 10318 12588 10324 12640
rect 10376 12628 10382 12640
rect 10413 12631 10471 12637
rect 10413 12628 10425 12631
rect 10376 12600 10425 12628
rect 10376 12588 10382 12600
rect 10413 12597 10425 12600
rect 10459 12597 10471 12631
rect 10413 12591 10471 12597
rect 12069 12631 12127 12637
rect 12069 12597 12081 12631
rect 12115 12628 12127 12631
rect 12434 12628 12440 12640
rect 12115 12600 12440 12628
rect 12115 12597 12127 12600
rect 12069 12591 12127 12597
rect 12434 12588 12440 12600
rect 12492 12588 12498 12640
rect 1104 12538 13708 12560
rect 1104 12486 2525 12538
rect 2577 12486 2589 12538
rect 2641 12486 2653 12538
rect 2705 12486 2717 12538
rect 2769 12486 2781 12538
rect 2833 12486 5676 12538
rect 5728 12486 5740 12538
rect 5792 12486 5804 12538
rect 5856 12486 5868 12538
rect 5920 12486 5932 12538
rect 5984 12486 8827 12538
rect 8879 12486 8891 12538
rect 8943 12486 8955 12538
rect 9007 12486 9019 12538
rect 9071 12486 9083 12538
rect 9135 12486 11978 12538
rect 12030 12486 12042 12538
rect 12094 12486 12106 12538
rect 12158 12486 12170 12538
rect 12222 12486 12234 12538
rect 12286 12486 13708 12538
rect 1104 12464 13708 12486
rect 4338 12384 4344 12436
rect 4396 12384 4402 12436
rect 4706 12384 4712 12436
rect 4764 12424 4770 12436
rect 4801 12427 4859 12433
rect 4801 12424 4813 12427
rect 4764 12396 4813 12424
rect 4764 12384 4770 12396
rect 4801 12393 4813 12396
rect 4847 12393 4859 12427
rect 4801 12387 4859 12393
rect 6178 12384 6184 12436
rect 6236 12424 6242 12436
rect 6273 12427 6331 12433
rect 6273 12424 6285 12427
rect 6236 12396 6285 12424
rect 6236 12384 6242 12396
rect 6273 12393 6285 12396
rect 6319 12393 6331 12427
rect 6273 12387 6331 12393
rect 6457 12427 6515 12433
rect 6457 12393 6469 12427
rect 6503 12424 6515 12427
rect 6730 12424 6736 12436
rect 6503 12396 6736 12424
rect 6503 12393 6515 12396
rect 6457 12387 6515 12393
rect 6730 12384 6736 12396
rect 6788 12384 6794 12436
rect 8202 12384 8208 12436
rect 8260 12384 8266 12436
rect 4614 12356 4620 12368
rect 4264 12328 4620 12356
rect 4264 12229 4292 12328
rect 4614 12316 4620 12328
rect 4672 12356 4678 12368
rect 5442 12356 5448 12368
rect 4672 12328 5448 12356
rect 4672 12316 4678 12328
rect 5442 12316 5448 12328
rect 5500 12356 5506 12368
rect 5500 12328 6224 12356
rect 5500 12316 5506 12328
rect 5537 12291 5595 12297
rect 5537 12288 5549 12291
rect 5276 12260 5549 12288
rect 4249 12223 4307 12229
rect 4249 12189 4261 12223
rect 4295 12189 4307 12223
rect 4249 12183 4307 12189
rect 4433 12223 4491 12229
rect 4433 12189 4445 12223
rect 4479 12189 4491 12223
rect 4433 12183 4491 12189
rect 4448 12152 4476 12183
rect 5074 12180 5080 12232
rect 5132 12180 5138 12232
rect 5166 12180 5172 12232
rect 5224 12180 5230 12232
rect 5276 12229 5304 12260
rect 5537 12257 5549 12260
rect 5583 12257 5595 12291
rect 6086 12288 6092 12300
rect 5537 12251 5595 12257
rect 5736 12260 6092 12288
rect 5261 12223 5319 12229
rect 5261 12189 5273 12223
rect 5307 12189 5319 12223
rect 5261 12183 5319 12189
rect 5442 12180 5448 12232
rect 5500 12180 5506 12232
rect 5736 12229 5764 12260
rect 6086 12248 6092 12260
rect 6144 12248 6150 12300
rect 5721 12223 5779 12229
rect 5721 12189 5733 12223
rect 5767 12189 5779 12223
rect 5721 12183 5779 12189
rect 5997 12223 6055 12229
rect 5997 12189 6009 12223
rect 6043 12220 6055 12223
rect 6196 12220 6224 12328
rect 7926 12248 7932 12300
rect 7984 12288 7990 12300
rect 9309 12291 9367 12297
rect 9309 12288 9321 12291
rect 7984 12260 9321 12288
rect 7984 12248 7990 12260
rect 9309 12257 9321 12260
rect 9355 12288 9367 12291
rect 10226 12288 10232 12300
rect 9355 12260 10232 12288
rect 9355 12257 9367 12260
rect 9309 12251 9367 12257
rect 10226 12248 10232 12260
rect 10284 12288 10290 12300
rect 11149 12291 11207 12297
rect 11149 12288 11161 12291
rect 10284 12260 11161 12288
rect 10284 12248 10290 12260
rect 11149 12257 11161 12260
rect 11195 12288 11207 12291
rect 11514 12288 11520 12300
rect 11195 12260 11520 12288
rect 11195 12257 11207 12260
rect 11149 12251 11207 12257
rect 11514 12248 11520 12260
rect 11572 12248 11578 12300
rect 6043 12192 6224 12220
rect 6043 12189 6055 12192
rect 5997 12183 6055 12189
rect 8386 12180 8392 12232
rect 8444 12180 8450 12232
rect 8570 12180 8576 12232
rect 8628 12220 8634 12232
rect 8665 12223 8723 12229
rect 8665 12220 8677 12223
rect 8628 12192 8677 12220
rect 8628 12180 8634 12192
rect 8665 12189 8677 12192
rect 8711 12189 8723 12223
rect 8665 12183 8723 12189
rect 5902 12152 5908 12164
rect 4448 12124 5908 12152
rect 5902 12112 5908 12124
rect 5960 12112 5966 12164
rect 6089 12155 6147 12161
rect 6089 12121 6101 12155
rect 6135 12121 6147 12155
rect 6089 12115 6147 12121
rect 6305 12155 6363 12161
rect 6305 12121 6317 12155
rect 6351 12152 6363 12155
rect 6914 12152 6920 12164
rect 6351 12124 6920 12152
rect 6351 12121 6363 12124
rect 6305 12115 6363 12121
rect 4154 12044 4160 12096
rect 4212 12084 4218 12096
rect 4522 12084 4528 12096
rect 4212 12056 4528 12084
rect 4212 12044 4218 12056
rect 4522 12044 4528 12056
rect 4580 12084 4586 12096
rect 6104 12084 6132 12115
rect 6914 12112 6920 12124
rect 6972 12112 6978 12164
rect 9585 12155 9643 12161
rect 9585 12121 9597 12155
rect 9631 12152 9643 12155
rect 9858 12152 9864 12164
rect 9631 12124 9864 12152
rect 9631 12121 9643 12124
rect 9585 12115 9643 12121
rect 9858 12112 9864 12124
rect 9916 12112 9922 12164
rect 10318 12112 10324 12164
rect 10376 12112 10382 12164
rect 11422 12112 11428 12164
rect 11480 12112 11486 12164
rect 12434 12112 12440 12164
rect 12492 12112 12498 12164
rect 6178 12084 6184 12096
rect 4580 12056 6184 12084
rect 4580 12044 4586 12056
rect 6178 12044 6184 12056
rect 6236 12084 6242 12096
rect 7190 12084 7196 12096
rect 6236 12056 7196 12084
rect 6236 12044 6242 12056
rect 7190 12044 7196 12056
rect 7248 12044 7254 12096
rect 8573 12087 8631 12093
rect 8573 12053 8585 12087
rect 8619 12084 8631 12087
rect 9398 12084 9404 12096
rect 8619 12056 9404 12084
rect 8619 12053 8631 12056
rect 8573 12047 8631 12053
rect 9398 12044 9404 12056
rect 9456 12044 9462 12096
rect 10870 12044 10876 12096
rect 10928 12084 10934 12096
rect 11057 12087 11115 12093
rect 11057 12084 11069 12087
rect 10928 12056 11069 12084
rect 10928 12044 10934 12056
rect 11057 12053 11069 12056
rect 11103 12053 11115 12087
rect 11057 12047 11115 12053
rect 12897 12087 12955 12093
rect 12897 12053 12909 12087
rect 12943 12084 12955 12087
rect 12986 12084 12992 12096
rect 12943 12056 12992 12084
rect 12943 12053 12955 12056
rect 12897 12047 12955 12053
rect 12986 12044 12992 12056
rect 13044 12044 13050 12096
rect 1104 11994 13708 12016
rect 1104 11942 3185 11994
rect 3237 11942 3249 11994
rect 3301 11942 3313 11994
rect 3365 11942 3377 11994
rect 3429 11942 3441 11994
rect 3493 11942 6336 11994
rect 6388 11942 6400 11994
rect 6452 11942 6464 11994
rect 6516 11942 6528 11994
rect 6580 11942 6592 11994
rect 6644 11942 9487 11994
rect 9539 11942 9551 11994
rect 9603 11942 9615 11994
rect 9667 11942 9679 11994
rect 9731 11942 9743 11994
rect 9795 11942 12638 11994
rect 12690 11942 12702 11994
rect 12754 11942 12766 11994
rect 12818 11942 12830 11994
rect 12882 11942 12894 11994
rect 12946 11942 13708 11994
rect 1104 11920 13708 11942
rect 1670 11840 1676 11892
rect 1728 11880 1734 11892
rect 4246 11880 4252 11892
rect 1728 11852 4252 11880
rect 1728 11840 1734 11852
rect 4246 11840 4252 11852
rect 4304 11840 4310 11892
rect 10226 11840 10232 11892
rect 10284 11840 10290 11892
rect 10778 11840 10784 11892
rect 10836 11880 10842 11892
rect 10836 11852 11284 11880
rect 10836 11840 10842 11852
rect 3605 11815 3663 11821
rect 3605 11812 3617 11815
rect 3174 11784 3617 11812
rect 3605 11781 3617 11784
rect 3651 11781 3663 11815
rect 3605 11775 3663 11781
rect 5166 11772 5172 11824
rect 5224 11812 5230 11824
rect 5965 11815 6023 11821
rect 5965 11812 5977 11815
rect 5224 11784 5977 11812
rect 5224 11772 5230 11784
rect 5965 11781 5977 11784
rect 6011 11781 6023 11815
rect 5965 11775 6023 11781
rect 6178 11772 6184 11824
rect 6236 11772 6242 11824
rect 8294 11812 8300 11824
rect 6288 11784 8300 11812
rect 3694 11704 3700 11756
rect 3752 11704 3758 11756
rect 5721 11747 5779 11753
rect 5721 11713 5733 11747
rect 5767 11744 5779 11747
rect 6288 11744 6316 11784
rect 8294 11772 8300 11784
rect 8352 11812 8358 11824
rect 8941 11815 8999 11821
rect 8941 11812 8953 11815
rect 8352 11784 8953 11812
rect 8352 11772 8358 11784
rect 8941 11781 8953 11784
rect 8987 11781 8999 11815
rect 8941 11775 8999 11781
rect 10962 11772 10968 11824
rect 11020 11772 11026 11824
rect 5767 11716 6316 11744
rect 6365 11747 6423 11753
rect 5767 11713 5779 11716
rect 5721 11707 5779 11713
rect 6365 11713 6377 11747
rect 6411 11713 6423 11747
rect 6365 11707 6423 11713
rect 1670 11636 1676 11688
rect 1728 11636 1734 11688
rect 1946 11636 1952 11688
rect 2004 11636 2010 11688
rect 5534 11636 5540 11688
rect 5592 11676 5598 11688
rect 6380 11676 6408 11707
rect 6546 11704 6552 11756
rect 6604 11704 6610 11756
rect 7009 11747 7067 11753
rect 7009 11744 7021 11747
rect 6932 11716 7021 11744
rect 5592 11648 6408 11676
rect 5592 11636 5598 11648
rect 3694 11568 3700 11620
rect 3752 11608 3758 11620
rect 6932 11608 6960 11716
rect 7009 11713 7021 11716
rect 7055 11744 7067 11747
rect 7098 11744 7104 11756
rect 7055 11716 7104 11744
rect 7055 11713 7067 11716
rect 7009 11707 7067 11713
rect 7098 11704 7104 11716
rect 7156 11704 7162 11756
rect 10873 11747 10931 11753
rect 10873 11713 10885 11747
rect 10919 11744 10931 11747
rect 10980 11744 11008 11772
rect 10919 11716 11008 11744
rect 10919 11713 10931 11716
rect 10873 11707 10931 11713
rect 11054 11704 11060 11756
rect 11112 11704 11118 11756
rect 11256 11744 11284 11852
rect 11422 11840 11428 11892
rect 11480 11880 11486 11892
rect 12161 11883 12219 11889
rect 12161 11880 12173 11883
rect 11480 11852 12173 11880
rect 11480 11840 11486 11852
rect 12161 11849 12173 11852
rect 12207 11849 12219 11883
rect 12161 11843 12219 11849
rect 11517 11747 11575 11753
rect 11517 11744 11529 11747
rect 11256 11716 11529 11744
rect 11517 11713 11529 11716
rect 11563 11713 11575 11747
rect 11517 11707 11575 11713
rect 11698 11704 11704 11756
rect 11756 11704 11762 11756
rect 11793 11747 11851 11753
rect 11793 11713 11805 11747
rect 11839 11713 11851 11747
rect 11793 11707 11851 11713
rect 11885 11747 11943 11753
rect 11885 11713 11897 11747
rect 11931 11744 11943 11747
rect 12342 11744 12348 11756
rect 11931 11716 12348 11744
rect 11931 11713 11943 11716
rect 11885 11707 11943 11713
rect 10594 11636 10600 11688
rect 10652 11676 10658 11688
rect 10965 11679 11023 11685
rect 10965 11676 10977 11679
rect 10652 11648 10977 11676
rect 10652 11636 10658 11648
rect 10965 11645 10977 11648
rect 11011 11676 11023 11679
rect 11808 11676 11836 11707
rect 12342 11704 12348 11716
rect 12400 11704 12406 11756
rect 11011 11648 11836 11676
rect 11011 11645 11023 11648
rect 10965 11639 11023 11645
rect 3752 11580 6960 11608
rect 3752 11568 3758 11580
rect 3421 11543 3479 11549
rect 3421 11509 3433 11543
rect 3467 11540 3479 11543
rect 3786 11540 3792 11552
rect 3467 11512 3792 11540
rect 3467 11509 3479 11512
rect 3421 11503 3479 11509
rect 3786 11500 3792 11512
rect 3844 11500 3850 11552
rect 4246 11500 4252 11552
rect 4304 11500 4310 11552
rect 4890 11500 4896 11552
rect 4948 11540 4954 11552
rect 5813 11543 5871 11549
rect 5813 11540 5825 11543
rect 4948 11512 5825 11540
rect 4948 11500 4954 11512
rect 5813 11509 5825 11512
rect 5859 11509 5871 11543
rect 5813 11503 5871 11509
rect 5997 11543 6055 11549
rect 5997 11509 6009 11543
rect 6043 11540 6055 11543
rect 6733 11543 6791 11549
rect 6733 11540 6745 11543
rect 6043 11512 6745 11540
rect 6043 11509 6055 11512
rect 5997 11503 6055 11509
rect 6733 11509 6745 11512
rect 6779 11509 6791 11543
rect 6733 11503 6791 11509
rect 6914 11500 6920 11552
rect 6972 11500 6978 11552
rect 1104 11450 13708 11472
rect 1104 11398 2525 11450
rect 2577 11398 2589 11450
rect 2641 11398 2653 11450
rect 2705 11398 2717 11450
rect 2769 11398 2781 11450
rect 2833 11398 5676 11450
rect 5728 11398 5740 11450
rect 5792 11398 5804 11450
rect 5856 11398 5868 11450
rect 5920 11398 5932 11450
rect 5984 11398 8827 11450
rect 8879 11398 8891 11450
rect 8943 11398 8955 11450
rect 9007 11398 9019 11450
rect 9071 11398 9083 11450
rect 9135 11398 11978 11450
rect 12030 11398 12042 11450
rect 12094 11398 12106 11450
rect 12158 11398 12170 11450
rect 12222 11398 12234 11450
rect 12286 11398 13708 11450
rect 1104 11376 13708 11398
rect 1946 11296 1952 11348
rect 2004 11336 2010 11348
rect 2133 11339 2191 11345
rect 2133 11336 2145 11339
rect 2004 11308 2145 11336
rect 2004 11296 2010 11308
rect 2133 11305 2145 11308
rect 2179 11305 2191 11339
rect 2133 11299 2191 11305
rect 2593 11339 2651 11345
rect 2593 11305 2605 11339
rect 2639 11336 2651 11339
rect 3421 11339 3479 11345
rect 3421 11336 3433 11339
rect 2639 11308 3433 11336
rect 2639 11305 2651 11308
rect 2593 11299 2651 11305
rect 3421 11305 3433 11308
rect 3467 11305 3479 11339
rect 3421 11299 3479 11305
rect 4709 11339 4767 11345
rect 4709 11305 4721 11339
rect 4755 11336 4767 11339
rect 5166 11336 5172 11348
rect 4755 11308 5172 11336
rect 4755 11305 4767 11308
rect 4709 11299 4767 11305
rect 5166 11296 5172 11308
rect 5224 11296 5230 11348
rect 5902 11296 5908 11348
rect 5960 11336 5966 11348
rect 6546 11336 6552 11348
rect 5960 11308 6552 11336
rect 5960 11296 5966 11308
rect 6546 11296 6552 11308
rect 6604 11336 6610 11348
rect 6917 11339 6975 11345
rect 6917 11336 6929 11339
rect 6604 11308 6929 11336
rect 6604 11296 6610 11308
rect 6917 11305 6929 11308
rect 6963 11305 6975 11339
rect 6917 11299 6975 11305
rect 9398 11296 9404 11348
rect 9456 11336 9462 11348
rect 9677 11339 9735 11345
rect 9677 11336 9689 11339
rect 9456 11308 9689 11336
rect 9456 11296 9462 11308
rect 9677 11305 9689 11308
rect 9723 11305 9735 11339
rect 9677 11299 9735 11305
rect 9858 11296 9864 11348
rect 9916 11336 9922 11348
rect 10137 11339 10195 11345
rect 10137 11336 10149 11339
rect 9916 11308 10149 11336
rect 9916 11296 9922 11308
rect 10137 11305 10149 11308
rect 10183 11305 10195 11339
rect 10137 11299 10195 11305
rect 11698 11296 11704 11348
rect 11756 11336 11762 11348
rect 11793 11339 11851 11345
rect 11793 11336 11805 11339
rect 11756 11308 11805 11336
rect 11756 11296 11762 11308
rect 11793 11305 11805 11308
rect 11839 11305 11851 11339
rect 11793 11299 11851 11305
rect 12342 11296 12348 11348
rect 12400 11296 12406 11348
rect 2409 11271 2467 11277
rect 2409 11237 2421 11271
rect 2455 11237 2467 11271
rect 2409 11231 2467 11237
rect 5077 11271 5135 11277
rect 5077 11237 5089 11271
rect 5123 11237 5135 11271
rect 5077 11231 5135 11237
rect 2317 11135 2375 11141
rect 2317 11101 2329 11135
rect 2363 11132 2375 11135
rect 2424 11132 2452 11231
rect 5092 11200 5120 11231
rect 10962 11228 10968 11280
rect 11020 11268 11026 11280
rect 11057 11271 11115 11277
rect 11057 11268 11069 11271
rect 11020 11240 11069 11268
rect 11020 11228 11026 11240
rect 11057 11237 11069 11240
rect 11103 11268 11115 11271
rect 12250 11268 12256 11280
rect 11103 11240 11468 11268
rect 11103 11237 11115 11240
rect 11057 11231 11115 11237
rect 5445 11203 5503 11209
rect 5445 11200 5457 11203
rect 5092 11172 5457 11200
rect 5445 11169 5457 11172
rect 5491 11169 5503 11203
rect 10980 11200 11008 11228
rect 11440 11212 11468 11240
rect 11900 11240 12256 11268
rect 5445 11163 5503 11169
rect 10428 11172 11008 11200
rect 11333 11203 11391 11209
rect 2958 11132 2964 11144
rect 2363 11104 2452 11132
rect 2700 11104 2964 11132
rect 2363 11101 2375 11104
rect 2317 11095 2375 11101
rect 2577 11067 2635 11073
rect 2577 11033 2589 11067
rect 2623 11064 2635 11067
rect 2700 11064 2728 11104
rect 2958 11092 2964 11104
rect 3016 11092 3022 11144
rect 3237 11135 3295 11141
rect 3237 11101 3249 11135
rect 3283 11132 3295 11135
rect 3513 11135 3571 11141
rect 3513 11132 3525 11135
rect 3283 11104 3525 11132
rect 3283 11101 3295 11104
rect 3237 11095 3295 11101
rect 3513 11101 3525 11104
rect 3559 11132 3571 11135
rect 4154 11132 4160 11144
rect 3559 11104 4160 11132
rect 3559 11101 3571 11104
rect 3513 11095 3571 11101
rect 4154 11092 4160 11104
rect 4212 11092 4218 11144
rect 4614 11092 4620 11144
rect 4672 11141 4678 11144
rect 4672 11132 4683 11141
rect 4672 11104 4717 11132
rect 4672 11095 4683 11104
rect 4672 11092 4678 11095
rect 4890 11092 4896 11144
rect 4948 11092 4954 11144
rect 5166 11092 5172 11144
rect 5224 11092 5230 11144
rect 6914 11132 6920 11144
rect 6578 11104 6920 11132
rect 6914 11092 6920 11104
rect 6972 11092 6978 11144
rect 8202 11092 8208 11144
rect 8260 11132 8266 11144
rect 10428 11141 10456 11172
rect 11333 11169 11345 11203
rect 11379 11169 11391 11203
rect 11333 11163 11391 11169
rect 10413 11135 10471 11141
rect 8260 11104 9996 11132
rect 8260 11092 8266 11104
rect 2623 11036 2728 11064
rect 2777 11067 2835 11073
rect 2623 11033 2635 11036
rect 2577 11027 2635 11033
rect 2777 11033 2789 11067
rect 2823 11033 2835 11067
rect 2777 11027 2835 11033
rect 3053 11067 3111 11073
rect 3053 11033 3065 11067
rect 3099 11033 3111 11067
rect 3053 11027 3111 11033
rect 4065 11067 4123 11073
rect 4065 11033 4077 11067
rect 4111 11064 4123 11067
rect 4246 11064 4252 11076
rect 4111 11036 4252 11064
rect 4111 11033 4123 11036
rect 4065 11027 4123 11033
rect 2406 10956 2412 11008
rect 2464 10996 2470 11008
rect 2792 10996 2820 11027
rect 2464 10968 2820 10996
rect 2464 10956 2470 10968
rect 2866 10956 2872 11008
rect 2924 10956 2930 11008
rect 3068 10996 3096 11027
rect 4246 11024 4252 11036
rect 4304 11064 4310 11076
rect 5184 11064 5212 11092
rect 4304 11036 5212 11064
rect 4304 11024 4310 11036
rect 7926 11024 7932 11076
rect 7984 11064 7990 11076
rect 9033 11067 9091 11073
rect 9033 11064 9045 11067
rect 7984 11036 9045 11064
rect 7984 11024 7990 11036
rect 9033 11033 9045 11036
rect 9079 11033 9091 11067
rect 9033 11027 9091 11033
rect 9214 11024 9220 11076
rect 9272 11064 9278 11076
rect 9861 11067 9919 11073
rect 9861 11064 9873 11067
rect 9272 11036 9873 11064
rect 9272 11024 9278 11036
rect 9861 11033 9873 11036
rect 9907 11033 9919 11067
rect 9968 11064 9996 11104
rect 10413 11101 10425 11135
rect 10459 11101 10471 11135
rect 10413 11095 10471 11101
rect 10502 11092 10508 11144
rect 10560 11092 10566 11144
rect 10594 11092 10600 11144
rect 10652 11092 10658 11144
rect 10778 11092 10784 11144
rect 10836 11092 10842 11144
rect 10870 11092 10876 11144
rect 10928 11092 10934 11144
rect 11348 11132 11376 11163
rect 11422 11160 11428 11212
rect 11480 11160 11486 11212
rect 11606 11160 11612 11212
rect 11664 11200 11670 11212
rect 11664 11172 11708 11200
rect 11664 11160 11670 11172
rect 11527 11135 11585 11141
rect 11348 11104 11468 11132
rect 10520 11064 10548 11092
rect 11054 11064 11060 11076
rect 9968 11036 11060 11064
rect 9861 11027 9919 11033
rect 11054 11024 11060 11036
rect 11112 11024 11118 11076
rect 11440 11064 11468 11104
rect 11527 11101 11539 11135
rect 11573 11126 11585 11135
rect 11790 11132 11796 11144
rect 11716 11126 11796 11132
rect 11573 11104 11796 11126
rect 11573 11101 11744 11104
rect 11527 11098 11744 11101
rect 11527 11095 11585 11098
rect 11790 11092 11796 11104
rect 11848 11132 11854 11144
rect 11900 11141 11928 11240
rect 12250 11228 12256 11240
rect 12308 11228 12314 11280
rect 12066 11160 12072 11212
rect 12124 11200 12130 11212
rect 12986 11200 12992 11212
rect 12124 11172 12992 11200
rect 12124 11160 12130 11172
rect 11885 11135 11943 11141
rect 11885 11132 11897 11135
rect 11848 11104 11897 11132
rect 11848 11092 11854 11104
rect 11885 11101 11897 11104
rect 11931 11101 11943 11135
rect 11885 11095 11943 11101
rect 12250 11092 12256 11144
rect 12308 11092 12314 11144
rect 12452 11141 12480 11172
rect 12986 11160 12992 11172
rect 13044 11160 13050 11212
rect 12437 11135 12495 11141
rect 12437 11101 12449 11135
rect 12483 11101 12495 11135
rect 12437 11095 12495 11101
rect 12529 11135 12587 11141
rect 12529 11101 12541 11135
rect 12575 11101 12587 11135
rect 12529 11095 12587 11101
rect 11977 11067 12035 11073
rect 11977 11064 11989 11067
rect 11440 11036 11989 11064
rect 11977 11033 11989 11036
rect 12023 11064 12035 11067
rect 12066 11064 12072 11076
rect 12023 11036 12072 11064
rect 12023 11033 12035 11036
rect 11977 11027 12035 11033
rect 12066 11024 12072 11036
rect 12124 11024 12130 11076
rect 12161 11067 12219 11073
rect 12161 11033 12173 11067
rect 12207 11064 12219 11067
rect 12342 11064 12348 11076
rect 12207 11036 12348 11064
rect 12207 11033 12219 11036
rect 12161 11027 12219 11033
rect 12342 11024 12348 11036
rect 12400 11024 12406 11076
rect 12544 11064 12572 11095
rect 12452 11036 12572 11064
rect 4522 10996 4528 11008
rect 3068 10968 4528 10996
rect 4522 10956 4528 10968
rect 4580 10956 4586 11008
rect 4614 10956 4620 11008
rect 4672 10996 4678 11008
rect 5442 10996 5448 11008
rect 4672 10968 5448 10996
rect 4672 10956 4678 10968
rect 5442 10956 5448 10968
rect 5500 10956 5506 11008
rect 8386 10956 8392 11008
rect 8444 10996 8450 11008
rect 9493 10999 9551 11005
rect 9493 10996 9505 10999
rect 8444 10968 9505 10996
rect 8444 10956 8450 10968
rect 9493 10965 9505 10968
rect 9539 10965 9551 10999
rect 9493 10959 9551 10965
rect 9661 10999 9719 11005
rect 9661 10965 9673 10999
rect 9707 10996 9719 10999
rect 9950 10996 9956 11008
rect 9707 10968 9956 10996
rect 9707 10965 9719 10968
rect 9661 10959 9719 10965
rect 9950 10956 9956 10968
rect 10008 10956 10014 11008
rect 11146 10956 11152 11008
rect 11204 10996 11210 11008
rect 11885 10999 11943 11005
rect 11885 10996 11897 10999
rect 11204 10968 11897 10996
rect 11204 10956 11210 10968
rect 11885 10965 11897 10968
rect 11931 10965 11943 10999
rect 11885 10959 11943 10965
rect 12250 10956 12256 11008
rect 12308 10996 12314 11008
rect 12452 10996 12480 11036
rect 12308 10968 12480 10996
rect 12308 10956 12314 10968
rect 12526 10956 12532 11008
rect 12584 10996 12590 11008
rect 12621 10999 12679 11005
rect 12621 10996 12633 10999
rect 12584 10968 12633 10996
rect 12584 10956 12590 10968
rect 12621 10965 12633 10968
rect 12667 10965 12679 10999
rect 12621 10959 12679 10965
rect 1104 10906 13708 10928
rect 1104 10854 3185 10906
rect 3237 10854 3249 10906
rect 3301 10854 3313 10906
rect 3365 10854 3377 10906
rect 3429 10854 3441 10906
rect 3493 10854 6336 10906
rect 6388 10854 6400 10906
rect 6452 10854 6464 10906
rect 6516 10854 6528 10906
rect 6580 10854 6592 10906
rect 6644 10854 9487 10906
rect 9539 10854 9551 10906
rect 9603 10854 9615 10906
rect 9667 10854 9679 10906
rect 9731 10854 9743 10906
rect 9795 10854 12638 10906
rect 12690 10854 12702 10906
rect 12754 10854 12766 10906
rect 12818 10854 12830 10906
rect 12882 10854 12894 10906
rect 12946 10854 13708 10906
rect 1104 10832 13708 10854
rect 1673 10795 1731 10801
rect 1673 10761 1685 10795
rect 1719 10792 1731 10795
rect 1719 10764 2084 10792
rect 1719 10761 1731 10764
rect 1673 10755 1731 10761
rect 2056 10733 2084 10764
rect 4154 10752 4160 10804
rect 4212 10792 4218 10804
rect 4249 10795 4307 10801
rect 4249 10792 4261 10795
rect 4212 10764 4261 10792
rect 4212 10752 4218 10764
rect 4249 10761 4261 10764
rect 4295 10761 4307 10795
rect 4249 10755 4307 10761
rect 5077 10795 5135 10801
rect 5077 10761 5089 10795
rect 5123 10792 5135 10795
rect 5534 10792 5540 10804
rect 5123 10764 5540 10792
rect 5123 10761 5135 10764
rect 5077 10755 5135 10761
rect 2041 10727 2099 10733
rect 2041 10693 2053 10727
rect 2087 10693 2099 10727
rect 2041 10687 2099 10693
rect 3050 10684 3056 10736
rect 3108 10684 3114 10736
rect 3786 10684 3792 10736
rect 3844 10684 3850 10736
rect 4005 10727 4063 10733
rect 4005 10693 4017 10727
rect 4051 10724 4063 10727
rect 4051 10696 4200 10724
rect 4051 10693 4063 10696
rect 4005 10687 4063 10693
rect 4172 10668 4200 10696
rect 1486 10616 1492 10668
rect 1544 10616 1550 10668
rect 4154 10616 4160 10668
rect 4212 10656 4218 10668
rect 4433 10659 4491 10665
rect 4433 10656 4445 10659
rect 4212 10628 4445 10656
rect 4212 10616 4218 10628
rect 4433 10625 4445 10628
rect 4479 10625 4491 10659
rect 4433 10619 4491 10625
rect 4985 10659 5043 10665
rect 4985 10625 4997 10659
rect 5031 10656 5043 10659
rect 5092 10656 5120 10755
rect 5534 10752 5540 10764
rect 5592 10752 5598 10804
rect 7009 10795 7067 10801
rect 7009 10792 7021 10795
rect 5828 10764 7021 10792
rect 5689 10727 5747 10733
rect 5689 10724 5701 10727
rect 5276 10696 5701 10724
rect 5276 10668 5304 10696
rect 5689 10693 5701 10696
rect 5735 10724 5747 10727
rect 5828 10724 5856 10764
rect 7009 10761 7021 10764
rect 7055 10792 7067 10795
rect 7653 10795 7711 10801
rect 7653 10792 7665 10795
rect 7055 10764 7665 10792
rect 7055 10761 7067 10764
rect 7009 10755 7067 10761
rect 7653 10761 7665 10764
rect 7699 10761 7711 10795
rect 7653 10755 7711 10761
rect 7745 10795 7803 10801
rect 7745 10761 7757 10795
rect 7791 10792 7803 10795
rect 8386 10792 8392 10804
rect 7791 10764 8392 10792
rect 7791 10761 7803 10764
rect 7745 10755 7803 10761
rect 8386 10752 8392 10764
rect 8444 10752 8450 10804
rect 8573 10795 8631 10801
rect 8573 10761 8585 10795
rect 8619 10792 8631 10795
rect 9398 10792 9404 10804
rect 8619 10764 9404 10792
rect 8619 10761 8631 10764
rect 8573 10755 8631 10761
rect 9398 10752 9404 10764
rect 9456 10792 9462 10804
rect 9582 10792 9588 10804
rect 9456 10764 9588 10792
rect 9456 10752 9462 10764
rect 9582 10752 9588 10764
rect 9640 10752 9646 10804
rect 10870 10792 10876 10804
rect 10060 10764 10876 10792
rect 5735 10696 5856 10724
rect 5735 10693 5747 10696
rect 5689 10687 5747 10693
rect 5902 10684 5908 10736
rect 5960 10684 5966 10736
rect 6825 10727 6883 10733
rect 6825 10724 6837 10727
rect 6288 10696 6837 10724
rect 5031 10628 5120 10656
rect 5031 10625 5043 10628
rect 4985 10619 5043 10625
rect 5258 10616 5264 10668
rect 5316 10616 5322 10668
rect 5350 10616 5356 10668
rect 5408 10656 5414 10668
rect 6288 10656 6316 10696
rect 6825 10693 6837 10696
rect 6871 10693 6883 10727
rect 6825 10687 6883 10693
rect 9125 10727 9183 10733
rect 9125 10693 9137 10727
rect 9171 10724 9183 10727
rect 9674 10724 9680 10736
rect 9171 10696 9680 10724
rect 9171 10693 9183 10696
rect 9125 10687 9183 10693
rect 5408 10628 6316 10656
rect 6549 10659 6607 10665
rect 5408 10616 5414 10628
rect 6549 10625 6561 10659
rect 6595 10656 6607 10659
rect 6730 10656 6736 10668
rect 6595 10628 6736 10656
rect 6595 10625 6607 10628
rect 6549 10619 6607 10625
rect 6730 10616 6736 10628
rect 6788 10616 6794 10668
rect 6840 10656 6868 10687
rect 9674 10684 9680 10696
rect 9732 10724 9738 10736
rect 10060 10724 10088 10764
rect 10870 10752 10876 10764
rect 10928 10752 10934 10804
rect 11422 10752 11428 10804
rect 11480 10792 11486 10804
rect 11698 10792 11704 10804
rect 11480 10764 11704 10792
rect 11480 10752 11486 10764
rect 11698 10752 11704 10764
rect 11756 10752 11762 10804
rect 9732 10696 10088 10724
rect 9732 10684 9738 10696
rect 10594 10684 10600 10736
rect 10652 10724 10658 10736
rect 10652 10696 11008 10724
rect 10652 10684 10658 10696
rect 7377 10659 7435 10665
rect 7377 10656 7389 10659
rect 6840 10628 7389 10656
rect 7377 10625 7389 10628
rect 7423 10625 7435 10659
rect 7377 10619 7435 10625
rect 7561 10659 7619 10665
rect 7561 10625 7573 10659
rect 7607 10625 7619 10659
rect 7561 10619 7619 10625
rect 7929 10659 7987 10665
rect 7929 10625 7941 10659
rect 7975 10656 7987 10659
rect 8021 10659 8079 10665
rect 8021 10656 8033 10659
rect 7975 10628 8033 10656
rect 7975 10625 7987 10628
rect 7929 10619 7987 10625
rect 8021 10625 8033 10628
rect 8067 10625 8079 10659
rect 8021 10619 8079 10625
rect 1670 10548 1676 10600
rect 1728 10588 1734 10600
rect 1765 10591 1823 10597
rect 1765 10588 1777 10591
rect 1728 10560 1777 10588
rect 1728 10548 1734 10560
rect 1765 10557 1777 10560
rect 1811 10557 1823 10591
rect 4522 10588 4528 10600
rect 1765 10551 1823 10557
rect 4080 10560 4528 10588
rect 3418 10412 3424 10464
rect 3476 10452 3482 10464
rect 3513 10455 3571 10461
rect 3513 10452 3525 10455
rect 3476 10424 3525 10452
rect 3476 10412 3482 10424
rect 3513 10421 3525 10424
rect 3559 10452 3571 10455
rect 3973 10455 4031 10461
rect 3973 10452 3985 10455
rect 3559 10424 3985 10452
rect 3559 10421 3571 10424
rect 3513 10415 3571 10421
rect 3973 10421 3985 10424
rect 4019 10452 4031 10455
rect 4080 10452 4108 10560
rect 4522 10548 4528 10560
rect 4580 10548 4586 10600
rect 4617 10591 4675 10597
rect 4617 10557 4629 10591
rect 4663 10588 4675 10591
rect 4798 10588 4804 10600
rect 4663 10560 4804 10588
rect 4663 10557 4675 10560
rect 4617 10551 4675 10557
rect 4798 10548 4804 10560
rect 4856 10548 4862 10600
rect 5902 10548 5908 10600
rect 5960 10588 5966 10600
rect 6365 10591 6423 10597
rect 6365 10588 6377 10591
rect 5960 10560 6377 10588
rect 5960 10548 5966 10560
rect 6365 10557 6377 10560
rect 6411 10588 6423 10591
rect 6822 10588 6828 10600
rect 6411 10560 6828 10588
rect 6411 10557 6423 10560
rect 6365 10551 6423 10557
rect 6822 10548 6828 10560
rect 6880 10548 6886 10600
rect 7576 10588 7604 10619
rect 8110 10616 8116 10668
rect 8168 10656 8174 10668
rect 8570 10656 8576 10668
rect 8168 10628 8576 10656
rect 8168 10616 8174 10628
rect 8570 10616 8576 10628
rect 8628 10656 8634 10668
rect 9306 10656 9312 10668
rect 8628 10628 9312 10656
rect 8628 10616 8634 10628
rect 9306 10616 9312 10628
rect 9364 10616 9370 10668
rect 9950 10656 9956 10668
rect 9416 10628 9956 10656
rect 7024 10560 7604 10588
rect 8665 10591 8723 10597
rect 4157 10523 4215 10529
rect 4157 10489 4169 10523
rect 4203 10520 4215 10523
rect 4430 10520 4436 10532
rect 4203 10492 4436 10520
rect 4203 10489 4215 10492
rect 4157 10483 4215 10489
rect 4430 10480 4436 10492
rect 4488 10480 4494 10532
rect 4706 10480 4712 10532
rect 4764 10520 4770 10532
rect 4764 10492 5212 10520
rect 4764 10480 4770 10492
rect 4019 10424 4108 10452
rect 4019 10421 4031 10424
rect 3973 10415 4031 10421
rect 4338 10412 4344 10464
rect 4396 10452 4402 10464
rect 4893 10455 4951 10461
rect 4893 10452 4905 10455
rect 4396 10424 4905 10452
rect 4396 10412 4402 10424
rect 4893 10421 4905 10424
rect 4939 10421 4951 10455
rect 5184 10452 5212 10492
rect 5350 10480 5356 10532
rect 5408 10520 5414 10532
rect 6733 10523 6791 10529
rect 5408 10492 5764 10520
rect 5408 10480 5414 10492
rect 5736 10461 5764 10492
rect 6733 10489 6745 10523
rect 6779 10520 6791 10523
rect 7024 10520 7052 10560
rect 8665 10557 8677 10591
rect 8711 10588 8723 10591
rect 9416 10588 9444 10628
rect 8711 10560 9444 10588
rect 8711 10557 8723 10560
rect 8665 10551 8723 10557
rect 9490 10548 9496 10600
rect 9548 10548 9554 10600
rect 9582 10548 9588 10600
rect 9640 10548 9646 10600
rect 9784 10597 9812 10628
rect 9950 10616 9956 10628
rect 10008 10616 10014 10668
rect 10318 10616 10324 10668
rect 10376 10656 10382 10668
rect 10689 10659 10747 10665
rect 10689 10656 10701 10659
rect 10376 10628 10701 10656
rect 10376 10616 10382 10628
rect 10689 10625 10701 10628
rect 10735 10656 10747 10659
rect 10778 10656 10784 10668
rect 10735 10628 10784 10656
rect 10735 10625 10747 10628
rect 10689 10619 10747 10625
rect 10778 10616 10784 10628
rect 10836 10616 10842 10668
rect 10980 10665 11008 10696
rect 12526 10684 12532 10736
rect 12584 10684 12590 10736
rect 10873 10659 10931 10665
rect 10873 10625 10885 10659
rect 10919 10625 10931 10659
rect 10873 10619 10931 10625
rect 10965 10659 11023 10665
rect 10965 10625 10977 10659
rect 11011 10625 11023 10659
rect 10965 10619 11023 10625
rect 11057 10659 11115 10665
rect 11057 10625 11069 10659
rect 11103 10656 11115 10659
rect 11146 10656 11152 10668
rect 11103 10628 11152 10656
rect 11103 10625 11115 10628
rect 11057 10619 11115 10625
rect 9677 10591 9735 10597
rect 9677 10557 9689 10591
rect 9723 10557 9735 10591
rect 9677 10551 9735 10557
rect 9769 10591 9827 10597
rect 9769 10557 9781 10591
rect 9815 10557 9827 10591
rect 10888 10588 10916 10619
rect 11146 10616 11152 10628
rect 11204 10616 11210 10668
rect 11514 10616 11520 10668
rect 11572 10616 11578 10668
rect 11238 10588 11244 10600
rect 10888 10560 11244 10588
rect 9769 10551 9827 10557
rect 6779 10492 7052 10520
rect 6779 10489 6791 10492
rect 6733 10483 6791 10489
rect 7024 10461 7052 10492
rect 7834 10480 7840 10532
rect 7892 10520 7898 10532
rect 8389 10523 8447 10529
rect 8389 10520 8401 10523
rect 7892 10492 8401 10520
rect 7892 10480 7898 10492
rect 8389 10489 8401 10492
rect 8435 10489 8447 10523
rect 8389 10483 8447 10489
rect 8478 10480 8484 10532
rect 8536 10520 8542 10532
rect 9125 10523 9183 10529
rect 9125 10520 9137 10523
rect 8536 10492 9137 10520
rect 8536 10480 8542 10492
rect 9125 10489 9137 10492
rect 9171 10520 9183 10523
rect 9214 10520 9220 10532
rect 9171 10492 9220 10520
rect 9171 10489 9183 10492
rect 9125 10483 9183 10489
rect 9214 10480 9220 10492
rect 9272 10520 9278 10532
rect 9272 10492 9444 10520
rect 9272 10480 9278 10492
rect 5537 10455 5595 10461
rect 5537 10452 5549 10455
rect 5184 10424 5549 10452
rect 4893 10415 4951 10421
rect 5537 10421 5549 10424
rect 5583 10421 5595 10455
rect 5537 10415 5595 10421
rect 5721 10455 5779 10461
rect 5721 10421 5733 10455
rect 5767 10421 5779 10455
rect 5721 10415 5779 10421
rect 7009 10455 7067 10461
rect 7009 10421 7021 10455
rect 7055 10421 7067 10455
rect 7009 10415 7067 10421
rect 7193 10455 7251 10461
rect 7193 10421 7205 10455
rect 7239 10452 7251 10455
rect 8110 10452 8116 10464
rect 7239 10424 8116 10452
rect 7239 10421 7251 10424
rect 7193 10415 7251 10421
rect 8110 10412 8116 10424
rect 8168 10412 8174 10464
rect 8202 10412 8208 10464
rect 8260 10412 8266 10464
rect 8570 10412 8576 10464
rect 8628 10452 8634 10464
rect 9309 10455 9367 10461
rect 9309 10452 9321 10455
rect 8628 10424 9321 10452
rect 8628 10412 8634 10424
rect 9309 10421 9321 10424
rect 9355 10421 9367 10455
rect 9416 10452 9444 10492
rect 9692 10452 9720 10551
rect 11238 10548 11244 10560
rect 11296 10548 11302 10600
rect 11333 10591 11391 10597
rect 11333 10557 11345 10591
rect 11379 10588 11391 10591
rect 11793 10591 11851 10597
rect 11793 10588 11805 10591
rect 11379 10560 11805 10588
rect 11379 10557 11391 10560
rect 11333 10551 11391 10557
rect 11793 10557 11805 10560
rect 11839 10557 11851 10591
rect 11793 10551 11851 10557
rect 9416 10424 9720 10452
rect 9309 10415 9367 10421
rect 11054 10412 11060 10464
rect 11112 10452 11118 10464
rect 12250 10452 12256 10464
rect 11112 10424 12256 10452
rect 11112 10412 11118 10424
rect 12250 10412 12256 10424
rect 12308 10412 12314 10464
rect 12342 10412 12348 10464
rect 12400 10452 12406 10464
rect 13265 10455 13323 10461
rect 13265 10452 13277 10455
rect 12400 10424 13277 10452
rect 12400 10412 12406 10424
rect 13265 10421 13277 10424
rect 13311 10421 13323 10455
rect 13265 10415 13323 10421
rect 1104 10362 13708 10384
rect 1104 10310 2525 10362
rect 2577 10310 2589 10362
rect 2641 10310 2653 10362
rect 2705 10310 2717 10362
rect 2769 10310 2781 10362
rect 2833 10310 5676 10362
rect 5728 10310 5740 10362
rect 5792 10310 5804 10362
rect 5856 10310 5868 10362
rect 5920 10310 5932 10362
rect 5984 10310 8827 10362
rect 8879 10310 8891 10362
rect 8943 10310 8955 10362
rect 9007 10310 9019 10362
rect 9071 10310 9083 10362
rect 9135 10310 11978 10362
rect 12030 10310 12042 10362
rect 12094 10310 12106 10362
rect 12158 10310 12170 10362
rect 12222 10310 12234 10362
rect 12286 10310 13708 10362
rect 1104 10288 13708 10310
rect 1486 10208 1492 10260
rect 1544 10248 1550 10260
rect 2317 10251 2375 10257
rect 2317 10248 2329 10251
rect 1544 10220 2329 10248
rect 1544 10208 1550 10220
rect 2317 10217 2329 10220
rect 2363 10217 2375 10251
rect 2317 10211 2375 10217
rect 2501 10251 2559 10257
rect 2501 10217 2513 10251
rect 2547 10217 2559 10251
rect 2501 10211 2559 10217
rect 2777 10251 2835 10257
rect 2777 10217 2789 10251
rect 2823 10248 2835 10251
rect 2958 10248 2964 10260
rect 2823 10220 2964 10248
rect 2823 10217 2835 10220
rect 2777 10211 2835 10217
rect 2516 10180 2544 10211
rect 2958 10208 2964 10220
rect 3016 10208 3022 10260
rect 3326 10208 3332 10260
rect 3384 10248 3390 10260
rect 3786 10248 3792 10260
rect 3384 10220 3792 10248
rect 3384 10208 3390 10220
rect 3786 10208 3792 10220
rect 3844 10248 3850 10260
rect 4706 10248 4712 10260
rect 3844 10220 4712 10248
rect 3844 10208 3850 10220
rect 4706 10208 4712 10220
rect 4764 10208 4770 10260
rect 6733 10251 6791 10257
rect 6733 10248 6745 10251
rect 4816 10220 6745 10248
rect 3881 10183 3939 10189
rect 3881 10180 3893 10183
rect 2516 10152 3893 10180
rect 3881 10149 3893 10152
rect 3927 10149 3939 10183
rect 3881 10143 3939 10149
rect 3605 10115 3663 10121
rect 3605 10081 3617 10115
rect 3651 10112 3663 10115
rect 4246 10112 4252 10124
rect 3651 10084 4252 10112
rect 3651 10081 3663 10084
rect 3605 10075 3663 10081
rect 2406 10004 2412 10056
rect 2464 10004 2470 10056
rect 2961 10047 3019 10053
rect 2961 10013 2973 10047
rect 3007 10044 3019 10047
rect 3326 10044 3332 10056
rect 3007 10016 3332 10044
rect 3007 10013 3019 10016
rect 2961 10007 3019 10013
rect 3326 10004 3332 10016
rect 3384 10004 3390 10056
rect 3418 10004 3424 10056
rect 3476 10004 3482 10056
rect 3988 10053 4016 10084
rect 4246 10072 4252 10084
rect 4304 10072 4310 10124
rect 3789 10047 3847 10053
rect 3789 10013 3801 10047
rect 3835 10013 3847 10047
rect 3789 10007 3847 10013
rect 3973 10047 4031 10053
rect 3973 10013 3985 10047
rect 4019 10013 4031 10047
rect 3973 10007 4031 10013
rect 4157 10047 4215 10053
rect 4157 10013 4169 10047
rect 4203 10044 4215 10047
rect 4203 10016 4292 10044
rect 4203 10013 4215 10016
rect 4157 10007 4215 10013
rect 2424 9976 2452 10004
rect 2685 9979 2743 9985
rect 2685 9976 2697 9979
rect 2424 9948 2697 9976
rect 2685 9945 2697 9948
rect 2731 9976 2743 9979
rect 3145 9979 3203 9985
rect 2731 9948 3096 9976
rect 2731 9945 2743 9948
rect 2685 9939 2743 9945
rect 2485 9911 2543 9917
rect 2485 9877 2497 9911
rect 2531 9908 2543 9911
rect 2866 9908 2872 9920
rect 2531 9880 2872 9908
rect 2531 9877 2543 9880
rect 2485 9871 2543 9877
rect 2866 9868 2872 9880
rect 2924 9868 2930 9920
rect 2958 9868 2964 9920
rect 3016 9908 3022 9920
rect 3068 9908 3096 9948
rect 3145 9945 3157 9979
rect 3191 9976 3203 9979
rect 3804 9976 3832 10007
rect 4264 9976 4292 10016
rect 4338 10004 4344 10056
rect 4396 10004 4402 10056
rect 4430 10004 4436 10056
rect 4488 10004 4494 10056
rect 4525 10047 4583 10053
rect 4525 10013 4537 10047
rect 4571 10044 4583 10047
rect 4816 10044 4844 10220
rect 6733 10217 6745 10220
rect 6779 10217 6791 10251
rect 6733 10211 6791 10217
rect 8205 10251 8263 10257
rect 8205 10217 8217 10251
rect 8251 10248 8263 10251
rect 9398 10248 9404 10260
rect 8251 10220 9404 10248
rect 8251 10217 8263 10220
rect 8205 10211 8263 10217
rect 9398 10208 9404 10220
rect 9456 10208 9462 10260
rect 11149 10251 11207 10257
rect 11149 10217 11161 10251
rect 11195 10217 11207 10251
rect 11149 10211 11207 10217
rect 8386 10140 8392 10192
rect 8444 10140 8450 10192
rect 9674 10180 9680 10192
rect 9324 10152 9680 10180
rect 4893 10115 4951 10121
rect 4893 10081 4905 10115
rect 4939 10112 4951 10115
rect 5166 10112 5172 10124
rect 4939 10084 5172 10112
rect 4939 10081 4951 10084
rect 4893 10075 4951 10081
rect 5166 10072 5172 10084
rect 5224 10072 5230 10124
rect 7377 10115 7435 10121
rect 7377 10081 7389 10115
rect 7423 10112 7435 10115
rect 8404 10112 8432 10140
rect 7423 10084 7696 10112
rect 7423 10081 7435 10084
rect 7377 10075 7435 10081
rect 4571 10016 4844 10044
rect 4571 10013 4583 10016
rect 4525 10007 4583 10013
rect 7098 10004 7104 10056
rect 7156 10044 7162 10056
rect 7469 10047 7527 10053
rect 7469 10044 7481 10047
rect 7156 10016 7481 10044
rect 7156 10004 7162 10016
rect 7469 10013 7481 10016
rect 7515 10013 7527 10047
rect 7469 10007 7527 10013
rect 4614 9976 4620 9988
rect 3191 9948 4200 9976
rect 4264 9948 4620 9976
rect 3191 9945 3203 9948
rect 3145 9939 3203 9945
rect 4172 9920 4200 9948
rect 4614 9936 4620 9948
rect 4672 9936 4678 9988
rect 4801 9979 4859 9985
rect 4801 9945 4813 9979
rect 4847 9976 4859 9979
rect 5169 9979 5227 9985
rect 5169 9976 5181 9979
rect 4847 9948 5181 9976
rect 4847 9945 4859 9948
rect 4801 9939 4859 9945
rect 5169 9945 5181 9948
rect 5215 9945 5227 9979
rect 7561 9979 7619 9985
rect 7561 9976 7573 9979
rect 6394 9948 7573 9976
rect 5169 9939 5227 9945
rect 7561 9945 7573 9948
rect 7607 9945 7619 9979
rect 7561 9939 7619 9945
rect 4062 9908 4068 9920
rect 3016 9880 4068 9908
rect 3016 9868 3022 9880
rect 4062 9868 4068 9880
rect 4120 9868 4126 9920
rect 4154 9868 4160 9920
rect 4212 9868 4218 9920
rect 5350 9868 5356 9920
rect 5408 9908 5414 9920
rect 6641 9911 6699 9917
rect 6641 9908 6653 9911
rect 5408 9880 6653 9908
rect 5408 9868 5414 9880
rect 6641 9877 6653 9880
rect 6687 9908 6699 9911
rect 7668 9908 7696 10084
rect 8128 10084 8432 10112
rect 8128 10053 8156 10084
rect 7837 10047 7895 10053
rect 7837 10013 7849 10047
rect 7883 10013 7895 10047
rect 7837 10007 7895 10013
rect 8113 10047 8171 10053
rect 8113 10013 8125 10047
rect 8159 10013 8171 10047
rect 8113 10007 8171 10013
rect 7852 9976 7880 10007
rect 8202 10004 8208 10056
rect 8260 10044 8266 10056
rect 8297 10047 8355 10053
rect 8297 10044 8309 10047
rect 8260 10016 8309 10044
rect 8260 10004 8266 10016
rect 8297 10013 8309 10016
rect 8343 10013 8355 10047
rect 8297 10007 8355 10013
rect 8478 10004 8484 10056
rect 8536 10004 8542 10056
rect 8573 10047 8631 10053
rect 8573 10013 8585 10047
rect 8619 10044 8631 10047
rect 8941 10047 8999 10053
rect 8941 10044 8953 10047
rect 8619 10016 8953 10044
rect 8619 10013 8631 10016
rect 8573 10007 8631 10013
rect 8941 10013 8953 10016
rect 8987 10013 8999 10047
rect 8941 10007 8999 10013
rect 9125 10047 9183 10053
rect 9125 10013 9137 10047
rect 9171 10044 9183 10047
rect 9324 10044 9352 10152
rect 9674 10140 9680 10152
rect 9732 10140 9738 10192
rect 11164 10180 11192 10211
rect 11238 10208 11244 10260
rect 11296 10248 11302 10260
rect 11425 10251 11483 10257
rect 11425 10248 11437 10251
rect 11296 10220 11437 10248
rect 11296 10208 11302 10220
rect 11425 10217 11437 10220
rect 11471 10217 11483 10251
rect 11425 10211 11483 10217
rect 11164 10152 11224 10180
rect 9950 10112 9956 10124
rect 9416 10084 9956 10112
rect 9416 10053 9444 10084
rect 9950 10072 9956 10084
rect 10008 10072 10014 10124
rect 11196 10112 11224 10152
rect 11790 10140 11796 10192
rect 11848 10180 11854 10192
rect 12713 10183 12771 10189
rect 12713 10180 12725 10183
rect 11848 10152 12725 10180
rect 11848 10140 11854 10152
rect 12713 10149 12725 10152
rect 12759 10149 12771 10183
rect 12713 10143 12771 10149
rect 11882 10112 11888 10124
rect 11196 10084 11888 10112
rect 11882 10072 11888 10084
rect 11940 10112 11946 10124
rect 11977 10115 12035 10121
rect 11977 10112 11989 10115
rect 11940 10084 11989 10112
rect 11940 10072 11946 10084
rect 11977 10081 11989 10084
rect 12023 10112 12035 10115
rect 12526 10112 12532 10124
rect 12023 10084 12532 10112
rect 12023 10081 12035 10084
rect 11977 10075 12035 10081
rect 12526 10072 12532 10084
rect 12584 10072 12590 10124
rect 9171 10016 9352 10044
rect 9401 10047 9459 10053
rect 9171 10013 9183 10016
rect 9125 10007 9183 10013
rect 9401 10013 9413 10047
rect 9447 10013 9459 10047
rect 9401 10007 9459 10013
rect 9677 10047 9735 10053
rect 9677 10013 9689 10047
rect 9723 10013 9735 10047
rect 11422 10044 11428 10056
rect 9677 10007 9735 10013
rect 10980 10016 11428 10044
rect 7852 9948 8340 9976
rect 6687 9880 7696 9908
rect 8021 9911 8079 9917
rect 6687 9877 6699 9880
rect 6641 9871 6699 9877
rect 8021 9877 8033 9911
rect 8067 9908 8079 9911
rect 8110 9908 8116 9920
rect 8067 9880 8116 9908
rect 8067 9877 8079 9880
rect 8021 9871 8079 9877
rect 8110 9868 8116 9880
rect 8168 9868 8174 9920
rect 8312 9908 8340 9948
rect 9214 9936 9220 9988
rect 9272 9976 9278 9988
rect 9585 9979 9643 9985
rect 9585 9976 9597 9979
rect 9272 9948 9597 9976
rect 9272 9936 9278 9948
rect 9585 9945 9597 9948
rect 9631 9945 9643 9979
rect 9585 9939 9643 9945
rect 8386 9908 8392 9920
rect 8312 9880 8392 9908
rect 8386 9868 8392 9880
rect 8444 9868 8450 9920
rect 8662 9868 8668 9920
rect 8720 9908 8726 9920
rect 8757 9911 8815 9917
rect 8757 9908 8769 9911
rect 8720 9880 8769 9908
rect 8720 9868 8726 9880
rect 8757 9877 8769 9880
rect 8803 9877 8815 9911
rect 8757 9871 8815 9877
rect 9306 9868 9312 9920
rect 9364 9868 9370 9920
rect 9692 9908 9720 10007
rect 10980 9985 11008 10016
rect 11422 10004 11428 10016
rect 11480 10004 11486 10056
rect 11609 10047 11667 10053
rect 11609 10013 11621 10047
rect 11655 10013 11667 10047
rect 11609 10007 11667 10013
rect 10965 9979 11023 9985
rect 10965 9945 10977 9979
rect 11011 9945 11023 9979
rect 10965 9939 11023 9945
rect 11181 9979 11239 9985
rect 11181 9945 11193 9979
rect 11227 9976 11239 9979
rect 11624 9976 11652 10007
rect 11698 10004 11704 10056
rect 11756 10004 11762 10056
rect 12066 10004 12072 10056
rect 12124 10004 12130 10056
rect 12345 10047 12403 10053
rect 12345 10013 12357 10047
rect 12391 10044 12403 10047
rect 13262 10044 13268 10056
rect 12391 10016 13268 10044
rect 12391 10013 12403 10016
rect 12345 10007 12403 10013
rect 13262 10004 13268 10016
rect 13320 10004 13326 10056
rect 11227 9948 12388 9976
rect 11227 9945 11239 9948
rect 11181 9939 11239 9945
rect 12360 9920 12388 9948
rect 12526 9936 12532 9988
rect 12584 9936 12590 9988
rect 10410 9908 10416 9920
rect 9692 9880 10416 9908
rect 10410 9868 10416 9880
rect 10468 9908 10474 9920
rect 11054 9908 11060 9920
rect 10468 9880 11060 9908
rect 10468 9868 10474 9880
rect 11054 9868 11060 9880
rect 11112 9868 11118 9920
rect 11330 9868 11336 9920
rect 11388 9868 11394 9920
rect 11422 9868 11428 9920
rect 11480 9908 11486 9920
rect 11790 9908 11796 9920
rect 11480 9880 11796 9908
rect 11480 9868 11486 9880
rect 11790 9868 11796 9880
rect 11848 9868 11854 9920
rect 11882 9868 11888 9920
rect 11940 9908 11946 9920
rect 12161 9911 12219 9917
rect 12161 9908 12173 9911
rect 11940 9880 12173 9908
rect 11940 9868 11946 9880
rect 12161 9877 12173 9880
rect 12207 9877 12219 9911
rect 12161 9871 12219 9877
rect 12342 9868 12348 9920
rect 12400 9908 12406 9920
rect 12437 9911 12495 9917
rect 12437 9908 12449 9911
rect 12400 9880 12449 9908
rect 12400 9868 12406 9880
rect 12437 9877 12449 9880
rect 12483 9877 12495 9911
rect 12437 9871 12495 9877
rect 1104 9818 13708 9840
rect 1104 9766 3185 9818
rect 3237 9766 3249 9818
rect 3301 9766 3313 9818
rect 3365 9766 3377 9818
rect 3429 9766 3441 9818
rect 3493 9766 6336 9818
rect 6388 9766 6400 9818
rect 6452 9766 6464 9818
rect 6516 9766 6528 9818
rect 6580 9766 6592 9818
rect 6644 9766 9487 9818
rect 9539 9766 9551 9818
rect 9603 9766 9615 9818
rect 9667 9766 9679 9818
rect 9731 9766 9743 9818
rect 9795 9766 12638 9818
rect 12690 9766 12702 9818
rect 12754 9766 12766 9818
rect 12818 9766 12830 9818
rect 12882 9766 12894 9818
rect 12946 9766 13708 9818
rect 1104 9744 13708 9766
rect 4709 9707 4767 9713
rect 4709 9673 4721 9707
rect 4755 9704 4767 9707
rect 5258 9704 5264 9716
rect 4755 9676 5264 9704
rect 4755 9673 4767 9676
rect 4709 9667 4767 9673
rect 5258 9664 5264 9676
rect 5316 9664 5322 9716
rect 8478 9664 8484 9716
rect 8536 9704 8542 9716
rect 9122 9704 9128 9716
rect 8536 9676 9128 9704
rect 8536 9664 8542 9676
rect 9122 9664 9128 9676
rect 9180 9664 9186 9716
rect 9677 9707 9735 9713
rect 9677 9673 9689 9707
rect 9723 9704 9735 9707
rect 9950 9704 9956 9716
rect 9723 9676 9956 9704
rect 9723 9673 9735 9676
rect 9677 9667 9735 9673
rect 9950 9664 9956 9676
rect 10008 9664 10014 9716
rect 10502 9664 10508 9716
rect 10560 9704 10566 9716
rect 11606 9704 11612 9716
rect 10560 9676 11612 9704
rect 10560 9664 10566 9676
rect 11606 9664 11612 9676
rect 11664 9704 11670 9716
rect 12066 9704 12072 9716
rect 11664 9676 12072 9704
rect 11664 9664 11670 9676
rect 12066 9664 12072 9676
rect 12124 9664 12130 9716
rect 2869 9639 2927 9645
rect 2869 9605 2881 9639
rect 2915 9636 2927 9639
rect 3050 9636 3056 9648
rect 2915 9608 3056 9636
rect 2915 9605 2927 9608
rect 2869 9599 2927 9605
rect 3050 9596 3056 9608
rect 3108 9596 3114 9648
rect 3694 9636 3700 9648
rect 3160 9608 3700 9636
rect 2961 9571 3019 9577
rect 2961 9537 2973 9571
rect 3007 9568 3019 9571
rect 3160 9568 3188 9608
rect 3694 9596 3700 9608
rect 3752 9596 3758 9648
rect 4246 9596 4252 9648
rect 4304 9636 4310 9648
rect 4525 9639 4583 9645
rect 4525 9636 4537 9639
rect 4304 9608 4537 9636
rect 4304 9596 4310 9608
rect 4525 9605 4537 9608
rect 4571 9605 4583 9639
rect 4525 9599 4583 9605
rect 4801 9639 4859 9645
rect 4801 9605 4813 9639
rect 4847 9636 4859 9639
rect 5350 9636 5356 9648
rect 4847 9608 5356 9636
rect 4847 9605 4859 9608
rect 4801 9599 4859 9605
rect 5350 9596 5356 9608
rect 5408 9596 5414 9648
rect 8110 9596 8116 9648
rect 8168 9636 8174 9648
rect 8205 9639 8263 9645
rect 8205 9636 8217 9639
rect 8168 9608 8217 9636
rect 8168 9596 8174 9608
rect 8205 9605 8217 9608
rect 8251 9605 8263 9639
rect 8205 9599 8263 9605
rect 9214 9596 9220 9648
rect 9272 9596 9278 9648
rect 12342 9596 12348 9648
rect 12400 9596 12406 9648
rect 3007 9540 3188 9568
rect 3237 9571 3295 9577
rect 3007 9537 3019 9540
rect 2961 9531 3019 9537
rect 3237 9537 3249 9571
rect 3283 9568 3295 9571
rect 4154 9568 4160 9580
rect 3283 9540 4160 9568
rect 3283 9537 3295 9540
rect 3237 9531 3295 9537
rect 2866 9460 2872 9512
rect 2924 9500 2930 9512
rect 2976 9500 3004 9531
rect 4154 9528 4160 9540
rect 4212 9528 4218 9580
rect 4338 9528 4344 9580
rect 4396 9528 4402 9580
rect 4430 9528 4436 9580
rect 4488 9528 4494 9580
rect 5077 9571 5135 9577
rect 5077 9537 5089 9571
rect 5123 9537 5135 9571
rect 5077 9531 5135 9537
rect 2924 9472 3004 9500
rect 2924 9460 2930 9472
rect 4522 9460 4528 9512
rect 4580 9500 4586 9512
rect 4893 9503 4951 9509
rect 4893 9500 4905 9503
rect 4580 9472 4905 9500
rect 4580 9460 4586 9472
rect 4893 9469 4905 9472
rect 4939 9469 4951 9503
rect 4893 9463 4951 9469
rect 3878 9392 3884 9444
rect 3936 9432 3942 9444
rect 4157 9435 4215 9441
rect 4157 9432 4169 9435
rect 3936 9404 4169 9432
rect 3936 9392 3942 9404
rect 4157 9401 4169 9404
rect 4203 9432 4215 9435
rect 5092 9432 5120 9531
rect 7926 9528 7932 9580
rect 7984 9528 7990 9580
rect 11514 9528 11520 9580
rect 11572 9528 11578 9580
rect 11054 9460 11060 9512
rect 11112 9500 11118 9512
rect 11793 9503 11851 9509
rect 11793 9500 11805 9503
rect 11112 9472 11805 9500
rect 11112 9460 11118 9472
rect 11793 9469 11805 9472
rect 11839 9469 11851 9503
rect 11793 9463 11851 9469
rect 13262 9460 13268 9512
rect 13320 9460 13326 9512
rect 4203 9404 5120 9432
rect 4203 9401 4215 9404
rect 4157 9395 4215 9401
rect 3142 9324 3148 9376
rect 3200 9324 3206 9376
rect 4798 9324 4804 9376
rect 4856 9324 4862 9376
rect 5261 9367 5319 9373
rect 5261 9333 5273 9367
rect 5307 9364 5319 9367
rect 5350 9364 5356 9376
rect 5307 9336 5356 9364
rect 5307 9333 5319 9336
rect 5261 9327 5319 9333
rect 5350 9324 5356 9336
rect 5408 9324 5414 9376
rect 1104 9274 13708 9296
rect 1104 9222 2525 9274
rect 2577 9222 2589 9274
rect 2641 9222 2653 9274
rect 2705 9222 2717 9274
rect 2769 9222 2781 9274
rect 2833 9222 5676 9274
rect 5728 9222 5740 9274
rect 5792 9222 5804 9274
rect 5856 9222 5868 9274
rect 5920 9222 5932 9274
rect 5984 9222 8827 9274
rect 8879 9222 8891 9274
rect 8943 9222 8955 9274
rect 9007 9222 9019 9274
rect 9071 9222 9083 9274
rect 9135 9222 11978 9274
rect 12030 9222 12042 9274
rect 12094 9222 12106 9274
rect 12158 9222 12170 9274
rect 12222 9222 12234 9274
rect 12286 9222 13708 9274
rect 1104 9200 13708 9222
rect 2777 9163 2835 9169
rect 2777 9129 2789 9163
rect 2823 9160 2835 9163
rect 3142 9160 3148 9172
rect 2823 9132 3148 9160
rect 2823 9129 2835 9132
rect 2777 9123 2835 9129
rect 3142 9120 3148 9132
rect 3200 9120 3206 9172
rect 4065 9163 4123 9169
rect 4065 9129 4077 9163
rect 4111 9129 4123 9163
rect 4065 9123 4123 9129
rect 4080 9092 4108 9123
rect 4154 9120 4160 9172
rect 4212 9160 4218 9172
rect 4249 9163 4307 9169
rect 4249 9160 4261 9163
rect 4212 9132 4261 9160
rect 4212 9120 4218 9132
rect 4249 9129 4261 9132
rect 4295 9129 4307 9163
rect 4249 9123 4307 9129
rect 8386 9120 8392 9172
rect 8444 9120 8450 9172
rect 8570 9120 8576 9172
rect 8628 9120 8634 9172
rect 11054 9120 11060 9172
rect 11112 9120 11118 9172
rect 12161 9163 12219 9169
rect 12161 9129 12173 9163
rect 12207 9160 12219 9163
rect 12342 9160 12348 9172
rect 12207 9132 12348 9160
rect 12207 9129 12219 9132
rect 12161 9123 12219 9129
rect 12342 9120 12348 9132
rect 12400 9120 12406 9172
rect 4338 9092 4344 9104
rect 4080 9064 4344 9092
rect 4338 9052 4344 9064
rect 4396 9092 4402 9104
rect 5442 9092 5448 9104
rect 4396 9064 5448 9092
rect 4396 9052 4402 9064
rect 5442 9052 5448 9064
rect 5500 9052 5506 9104
rect 11330 9052 11336 9104
rect 11388 9092 11394 9104
rect 11388 9064 11744 9092
rect 11388 9052 11394 9064
rect 6822 9024 6828 9036
rect 5276 8996 6828 9024
rect 5276 8965 5304 8996
rect 6822 8984 6828 8996
rect 6880 8984 6886 9036
rect 6914 8984 6920 9036
rect 6972 9024 6978 9036
rect 8202 9024 8208 9036
rect 6972 8996 8208 9024
rect 6972 8984 6978 8996
rect 8202 8984 8208 8996
rect 8260 8984 8266 9036
rect 11425 9027 11483 9033
rect 11425 9024 11437 9027
rect 10612 8996 11437 9024
rect 2409 8959 2467 8965
rect 2409 8925 2421 8959
rect 2455 8956 2467 8959
rect 5261 8959 5319 8965
rect 2455 8928 2636 8956
rect 2455 8925 2467 8928
rect 2409 8919 2467 8925
rect 1946 8780 1952 8832
rect 2004 8820 2010 8832
rect 2608 8829 2636 8928
rect 5261 8925 5273 8959
rect 5307 8925 5319 8959
rect 5261 8919 5319 8925
rect 5350 8916 5356 8968
rect 5408 8916 5414 8968
rect 5442 8916 5448 8968
rect 5500 8956 5506 8968
rect 5537 8959 5595 8965
rect 5537 8956 5549 8959
rect 5500 8928 5549 8956
rect 5500 8916 5506 8928
rect 5537 8925 5549 8928
rect 5583 8925 5595 8959
rect 5537 8919 5595 8925
rect 5629 8959 5687 8965
rect 5629 8925 5641 8959
rect 5675 8925 5687 8959
rect 5629 8919 5687 8925
rect 2958 8848 2964 8900
rect 3016 8848 3022 8900
rect 3878 8848 3884 8900
rect 3936 8848 3942 8900
rect 4097 8891 4155 8897
rect 4097 8857 4109 8891
rect 4143 8888 4155 8891
rect 4430 8888 4436 8900
rect 4143 8860 4436 8888
rect 4143 8857 4155 8860
rect 4097 8851 4155 8857
rect 4430 8848 4436 8860
rect 4488 8888 4494 8900
rect 5166 8888 5172 8900
rect 4488 8860 5172 8888
rect 4488 8848 4494 8860
rect 5166 8848 5172 8860
rect 5224 8888 5230 8900
rect 5644 8888 5672 8919
rect 6546 8916 6552 8968
rect 6604 8916 6610 8968
rect 8570 8916 8576 8968
rect 8628 8916 8634 8968
rect 10318 8916 10324 8968
rect 10376 8956 10382 8968
rect 10612 8965 10640 8996
rect 11425 8993 11437 8996
rect 11471 8993 11483 9027
rect 11425 8987 11483 8993
rect 11606 8984 11612 9036
rect 11664 8984 11670 9036
rect 11716 9033 11744 9064
rect 11701 9027 11759 9033
rect 11701 8993 11713 9027
rect 11747 8993 11759 9027
rect 11701 8987 11759 8993
rect 11885 9027 11943 9033
rect 11885 8993 11897 9027
rect 11931 9024 11943 9027
rect 12621 9027 12679 9033
rect 12621 9024 12633 9027
rect 11931 8996 12633 9024
rect 11931 8993 11943 8996
rect 11885 8987 11943 8993
rect 12621 8993 12633 8996
rect 12667 8993 12679 9027
rect 12621 8987 12679 8993
rect 13262 8984 13268 9036
rect 13320 8984 13326 9036
rect 10413 8959 10471 8965
rect 10413 8956 10425 8959
rect 10376 8928 10425 8956
rect 10376 8916 10382 8928
rect 10413 8925 10425 8928
rect 10459 8925 10471 8959
rect 10413 8919 10471 8925
rect 10597 8959 10655 8965
rect 10597 8925 10609 8959
rect 10643 8925 10655 8959
rect 10597 8919 10655 8925
rect 10689 8959 10747 8965
rect 10689 8925 10701 8959
rect 10735 8925 10747 8959
rect 10689 8919 10747 8925
rect 5224 8860 5672 8888
rect 8588 8888 8616 8916
rect 8757 8891 8815 8897
rect 8757 8888 8769 8891
rect 8588 8860 8769 8888
rect 5224 8848 5230 8860
rect 8757 8857 8769 8860
rect 8803 8857 8815 8891
rect 8757 8851 8815 8857
rect 9398 8848 9404 8900
rect 9456 8888 9462 8900
rect 10042 8888 10048 8900
rect 9456 8860 10048 8888
rect 9456 8848 9462 8860
rect 10042 8848 10048 8860
rect 10100 8888 10106 8900
rect 10704 8888 10732 8919
rect 10778 8916 10784 8968
rect 10836 8916 10842 8968
rect 11793 8959 11851 8965
rect 11793 8925 11805 8959
rect 11839 8925 11851 8959
rect 11793 8919 11851 8925
rect 12069 8959 12127 8965
rect 12069 8925 12081 8959
rect 12115 8956 12127 8959
rect 12342 8956 12348 8968
rect 12115 8928 12348 8956
rect 12115 8925 12127 8928
rect 12069 8919 12127 8925
rect 10100 8860 10732 8888
rect 10100 8848 10106 8860
rect 11698 8848 11704 8900
rect 11756 8888 11762 8900
rect 11808 8888 11836 8919
rect 12342 8916 12348 8928
rect 12400 8916 12406 8968
rect 11756 8860 11836 8888
rect 11756 8848 11762 8860
rect 2225 8823 2283 8829
rect 2225 8820 2237 8823
rect 2004 8792 2237 8820
rect 2004 8780 2010 8792
rect 2225 8789 2237 8792
rect 2271 8789 2283 8823
rect 2225 8783 2283 8789
rect 2593 8823 2651 8829
rect 2593 8789 2605 8823
rect 2639 8789 2651 8823
rect 2593 8783 2651 8789
rect 2761 8823 2819 8829
rect 2761 8789 2773 8823
rect 2807 8820 2819 8823
rect 3510 8820 3516 8832
rect 2807 8792 3516 8820
rect 2807 8789 2819 8792
rect 2761 8783 2819 8789
rect 3510 8780 3516 8792
rect 3568 8780 3574 8832
rect 5813 8823 5871 8829
rect 5813 8789 5825 8823
rect 5859 8820 5871 8823
rect 8386 8820 8392 8832
rect 5859 8792 8392 8820
rect 5859 8789 5871 8792
rect 5813 8783 5871 8789
rect 8386 8780 8392 8792
rect 8444 8780 8450 8832
rect 8557 8823 8615 8829
rect 8557 8789 8569 8823
rect 8603 8820 8615 8823
rect 9416 8820 9444 8848
rect 8603 8792 9444 8820
rect 8603 8789 8615 8792
rect 8557 8783 8615 8789
rect 1104 8730 13708 8752
rect 1104 8678 3185 8730
rect 3237 8678 3249 8730
rect 3301 8678 3313 8730
rect 3365 8678 3377 8730
rect 3429 8678 3441 8730
rect 3493 8678 6336 8730
rect 6388 8678 6400 8730
rect 6452 8678 6464 8730
rect 6516 8678 6528 8730
rect 6580 8678 6592 8730
rect 6644 8678 9487 8730
rect 9539 8678 9551 8730
rect 9603 8678 9615 8730
rect 9667 8678 9679 8730
rect 9731 8678 9743 8730
rect 9795 8678 12638 8730
rect 12690 8678 12702 8730
rect 12754 8678 12766 8730
rect 12818 8678 12830 8730
rect 12882 8678 12894 8730
rect 12946 8678 13708 8730
rect 1104 8656 13708 8678
rect 3421 8619 3479 8625
rect 3421 8585 3433 8619
rect 3467 8585 3479 8619
rect 3421 8579 3479 8585
rect 1946 8508 1952 8560
rect 2004 8508 2010 8560
rect 2958 8508 2964 8560
rect 3016 8508 3022 8560
rect 3436 8548 3464 8579
rect 3510 8576 3516 8628
rect 3568 8576 3574 8628
rect 3878 8616 3884 8628
rect 3712 8588 3884 8616
rect 3712 8557 3740 8588
rect 3878 8576 3884 8588
rect 3936 8576 3942 8628
rect 6730 8576 6736 8628
rect 6788 8616 6794 8628
rect 6788 8588 7420 8616
rect 6788 8576 6794 8588
rect 3697 8551 3755 8557
rect 3697 8548 3709 8551
rect 3436 8520 3709 8548
rect 3697 8517 3709 8520
rect 3743 8517 3755 8551
rect 7392 8548 7420 8588
rect 7650 8576 7656 8628
rect 7708 8576 7714 8628
rect 8294 8576 8300 8628
rect 8352 8616 8358 8628
rect 8478 8616 8484 8628
rect 8352 8588 8484 8616
rect 8352 8576 8358 8588
rect 8478 8576 8484 8588
rect 8536 8576 8542 8628
rect 8662 8576 8668 8628
rect 8720 8616 8726 8628
rect 8720 8588 8892 8616
rect 8720 8576 8726 8588
rect 7805 8551 7863 8557
rect 7805 8548 7817 8551
rect 3697 8511 3755 8517
rect 6748 8520 7328 8548
rect 7392 8520 7817 8548
rect 1670 8440 1676 8492
rect 1728 8440 1734 8492
rect 3881 8483 3939 8489
rect 3881 8449 3893 8483
rect 3927 8480 3939 8483
rect 4338 8480 4344 8492
rect 3927 8452 4344 8480
rect 3927 8449 3939 8452
rect 3881 8443 3939 8449
rect 4338 8440 4344 8452
rect 4396 8440 4402 8492
rect 5350 8440 5356 8492
rect 5408 8480 5414 8492
rect 6748 8489 6776 8520
rect 6733 8483 6791 8489
rect 6733 8480 6745 8483
rect 5408 8452 6745 8480
rect 5408 8440 5414 8452
rect 6733 8449 6745 8452
rect 6779 8449 6791 8483
rect 6733 8443 6791 8449
rect 6822 8440 6828 8492
rect 6880 8480 6886 8492
rect 7300 8489 7328 8520
rect 7805 8517 7817 8520
rect 7851 8517 7863 8551
rect 7805 8511 7863 8517
rect 7926 8508 7932 8560
rect 7984 8557 7990 8560
rect 8864 8557 8892 8588
rect 7984 8551 8033 8557
rect 7984 8517 7987 8551
rect 8021 8517 8033 8551
rect 7984 8511 8033 8517
rect 8849 8551 8907 8557
rect 8849 8517 8861 8551
rect 8895 8517 8907 8551
rect 8849 8511 8907 8517
rect 7984 8508 7990 8511
rect 9214 8508 9220 8560
rect 9272 8548 9278 8560
rect 10594 8548 10600 8560
rect 9272 8520 10600 8548
rect 9272 8508 9278 8520
rect 7101 8483 7159 8489
rect 7101 8480 7113 8483
rect 6880 8452 7113 8480
rect 6880 8440 6886 8452
rect 7101 8449 7113 8452
rect 7147 8449 7159 8483
rect 7101 8443 7159 8449
rect 7285 8483 7343 8489
rect 7285 8449 7297 8483
rect 7331 8449 7343 8483
rect 8113 8483 8171 8489
rect 8113 8480 8125 8483
rect 7285 8443 7343 8449
rect 7576 8452 8125 8480
rect 6638 8372 6644 8424
rect 6696 8372 6702 8424
rect 7009 8415 7067 8421
rect 7009 8381 7021 8415
rect 7055 8412 7067 8415
rect 7576 8412 7604 8452
rect 8113 8449 8125 8452
rect 8159 8449 8171 8483
rect 8113 8443 8171 8449
rect 8205 8483 8263 8489
rect 8205 8449 8217 8483
rect 8251 8449 8263 8483
rect 8205 8443 8263 8449
rect 7055 8384 7604 8412
rect 7055 8381 7067 8384
rect 7009 8375 7067 8381
rect 7834 8372 7840 8424
rect 7892 8412 7898 8424
rect 7892 8384 8064 8412
rect 7892 8372 7898 8384
rect 8036 8344 8064 8384
rect 8220 8344 8248 8443
rect 8386 8440 8392 8492
rect 8444 8480 8450 8492
rect 8573 8483 8631 8489
rect 8573 8480 8585 8483
rect 8444 8452 8585 8480
rect 8444 8440 8450 8452
rect 8573 8449 8585 8452
rect 8619 8449 8631 8483
rect 8573 8443 8631 8449
rect 8662 8440 8668 8492
rect 8720 8440 8726 8492
rect 10520 8489 10548 8520
rect 10594 8508 10600 8520
rect 10652 8548 10658 8560
rect 11330 8548 11336 8560
rect 10652 8520 11336 8548
rect 10652 8508 10658 8520
rect 11330 8508 11336 8520
rect 11388 8548 11394 8560
rect 11882 8548 11888 8560
rect 11388 8520 11888 8548
rect 11388 8508 11394 8520
rect 11882 8508 11888 8520
rect 11940 8508 11946 8560
rect 10505 8483 10563 8489
rect 10505 8449 10517 8483
rect 10551 8449 10563 8483
rect 10505 8443 10563 8449
rect 10689 8483 10747 8489
rect 10689 8449 10701 8483
rect 10735 8480 10747 8483
rect 10870 8480 10876 8492
rect 10735 8452 10876 8480
rect 10735 8449 10747 8452
rect 10689 8443 10747 8449
rect 10870 8440 10876 8452
rect 10928 8440 10934 8492
rect 8478 8372 8484 8424
rect 8536 8372 8542 8424
rect 8036 8316 8248 8344
rect 4706 8236 4712 8288
rect 4764 8276 4770 8288
rect 6730 8276 6736 8288
rect 4764 8248 6736 8276
rect 4764 8236 4770 8248
rect 6730 8236 6736 8248
rect 6788 8236 6794 8288
rect 7282 8236 7288 8288
rect 7340 8236 7346 8288
rect 7877 8279 7935 8285
rect 7877 8245 7889 8279
rect 7923 8276 7935 8279
rect 8036 8276 8064 8316
rect 8386 8304 8392 8356
rect 8444 8304 8450 8356
rect 7923 8248 8064 8276
rect 7923 8245 7935 8248
rect 7877 8239 7935 8245
rect 8662 8236 8668 8288
rect 8720 8276 8726 8288
rect 8849 8279 8907 8285
rect 8849 8276 8861 8279
rect 8720 8248 8861 8276
rect 8720 8236 8726 8248
rect 8849 8245 8861 8248
rect 8895 8245 8907 8279
rect 8849 8239 8907 8245
rect 10134 8236 10140 8288
rect 10192 8276 10198 8288
rect 10597 8279 10655 8285
rect 10597 8276 10609 8279
rect 10192 8248 10609 8276
rect 10192 8236 10198 8248
rect 10597 8245 10609 8248
rect 10643 8276 10655 8279
rect 10778 8276 10784 8288
rect 10643 8248 10784 8276
rect 10643 8245 10655 8248
rect 10597 8239 10655 8245
rect 10778 8236 10784 8248
rect 10836 8236 10842 8288
rect 1104 8186 13708 8208
rect 1104 8134 2525 8186
rect 2577 8134 2589 8186
rect 2641 8134 2653 8186
rect 2705 8134 2717 8186
rect 2769 8134 2781 8186
rect 2833 8134 5676 8186
rect 5728 8134 5740 8186
rect 5792 8134 5804 8186
rect 5856 8134 5868 8186
rect 5920 8134 5932 8186
rect 5984 8134 8827 8186
rect 8879 8134 8891 8186
rect 8943 8134 8955 8186
rect 9007 8134 9019 8186
rect 9071 8134 9083 8186
rect 9135 8134 11978 8186
rect 12030 8134 12042 8186
rect 12094 8134 12106 8186
rect 12158 8134 12170 8186
rect 12222 8134 12234 8186
rect 12286 8134 13708 8186
rect 1104 8112 13708 8134
rect 2777 8075 2835 8081
rect 2777 8041 2789 8075
rect 2823 8072 2835 8075
rect 2958 8072 2964 8084
rect 2823 8044 2964 8072
rect 2823 8041 2835 8044
rect 2777 8035 2835 8041
rect 2958 8032 2964 8044
rect 3016 8032 3022 8084
rect 4706 8032 4712 8084
rect 4764 8032 4770 8084
rect 4816 8044 5028 8072
rect 4338 7964 4344 8016
rect 4396 8004 4402 8016
rect 4816 8004 4844 8044
rect 5000 8013 5028 8044
rect 9692 8044 11008 8072
rect 4396 7976 4844 8004
rect 4893 8007 4951 8013
rect 4396 7964 4402 7976
rect 4893 7973 4905 8007
rect 4939 7973 4951 8007
rect 4893 7967 4951 7973
rect 4985 8007 5043 8013
rect 4985 7973 4997 8007
rect 5031 8004 5043 8007
rect 7929 8007 7987 8013
rect 7929 8004 7941 8007
rect 5031 7976 7941 8004
rect 5031 7973 5043 7976
rect 4985 7967 5043 7973
rect 7929 7973 7941 7976
rect 7975 8004 7987 8007
rect 8478 8004 8484 8016
rect 7975 7976 8484 8004
rect 7975 7973 7987 7976
rect 7929 7967 7987 7973
rect 4908 7936 4936 7967
rect 8478 7964 8484 7976
rect 8536 7964 8542 8016
rect 4908 7908 5488 7936
rect 2866 7828 2872 7880
rect 2924 7828 2930 7880
rect 5166 7828 5172 7880
rect 5224 7828 5230 7880
rect 5261 7871 5319 7877
rect 5261 7837 5273 7871
rect 5307 7868 5319 7871
rect 5350 7868 5356 7880
rect 5307 7840 5356 7868
rect 5307 7837 5319 7840
rect 5261 7831 5319 7837
rect 4430 7760 4436 7812
rect 4488 7800 4494 7812
rect 5276 7800 5304 7831
rect 5350 7828 5356 7840
rect 5408 7828 5414 7880
rect 5460 7877 5488 7908
rect 5445 7871 5503 7877
rect 5445 7837 5457 7871
rect 5491 7837 5503 7871
rect 5445 7831 5503 7837
rect 7650 7828 7656 7880
rect 7708 7868 7714 7880
rect 8113 7871 8171 7877
rect 8113 7868 8125 7871
rect 7708 7840 8125 7868
rect 7708 7828 7714 7840
rect 8113 7837 8125 7840
rect 8159 7837 8171 7871
rect 8113 7831 8171 7837
rect 8294 7828 8300 7880
rect 8352 7868 8358 7880
rect 8573 7871 8631 7877
rect 8573 7868 8585 7871
rect 8352 7840 8585 7868
rect 8352 7828 8358 7840
rect 8573 7837 8585 7840
rect 8619 7837 8631 7871
rect 8573 7831 8631 7837
rect 8754 7828 8760 7880
rect 8812 7828 8818 7880
rect 9692 7877 9720 8044
rect 10045 8007 10103 8013
rect 10045 7973 10057 8007
rect 10091 8004 10103 8007
rect 10134 8004 10140 8016
rect 10091 7976 10140 8004
rect 10091 7973 10103 7976
rect 10045 7967 10103 7973
rect 10134 7964 10140 7976
rect 10192 7964 10198 8016
rect 10505 7939 10563 7945
rect 10505 7936 10517 7939
rect 10244 7908 10517 7936
rect 9677 7871 9735 7877
rect 9677 7837 9689 7871
rect 9723 7837 9735 7871
rect 9677 7831 9735 7837
rect 9950 7828 9956 7880
rect 10008 7828 10014 7880
rect 10042 7828 10048 7880
rect 10100 7868 10106 7880
rect 10244 7877 10272 7908
rect 10505 7905 10517 7908
rect 10551 7905 10563 7939
rect 10505 7899 10563 7905
rect 10594 7896 10600 7948
rect 10652 7936 10658 7948
rect 10980 7945 11008 8044
rect 12342 8004 12348 8016
rect 11348 7976 12348 8004
rect 10781 7939 10839 7945
rect 10781 7936 10793 7939
rect 10652 7908 10793 7936
rect 10652 7896 10658 7908
rect 10781 7905 10793 7908
rect 10827 7905 10839 7939
rect 10781 7899 10839 7905
rect 10965 7939 11023 7945
rect 10965 7905 10977 7939
rect 11011 7936 11023 7939
rect 11146 7936 11152 7948
rect 11011 7908 11152 7936
rect 11011 7905 11023 7908
rect 10965 7899 11023 7905
rect 11146 7896 11152 7908
rect 11204 7896 11210 7948
rect 10137 7871 10195 7877
rect 10137 7868 10149 7871
rect 10100 7840 10149 7868
rect 10100 7828 10106 7840
rect 10137 7837 10149 7840
rect 10183 7837 10195 7871
rect 10137 7831 10195 7837
rect 10229 7871 10287 7877
rect 10229 7837 10241 7871
rect 10275 7837 10287 7871
rect 10229 7831 10287 7837
rect 10318 7828 10324 7880
rect 10376 7868 10382 7880
rect 10413 7871 10471 7877
rect 10413 7868 10425 7871
rect 10376 7840 10425 7868
rect 10376 7828 10382 7840
rect 10413 7837 10425 7840
rect 10459 7837 10471 7871
rect 10413 7831 10471 7837
rect 10689 7871 10747 7877
rect 10689 7837 10701 7871
rect 10735 7837 10747 7871
rect 10689 7831 10747 7837
rect 4488 7772 5304 7800
rect 8205 7803 8263 7809
rect 4488 7760 4494 7772
rect 8205 7769 8217 7803
rect 8251 7800 8263 7803
rect 8665 7803 8723 7809
rect 8665 7800 8677 7803
rect 8251 7772 8677 7800
rect 8251 7769 8263 7772
rect 8205 7763 8263 7769
rect 8665 7769 8677 7772
rect 8711 7769 8723 7803
rect 8665 7763 8723 7769
rect 9585 7803 9643 7809
rect 9585 7769 9597 7803
rect 9631 7800 9643 7803
rect 9968 7800 9996 7828
rect 9631 7772 9996 7800
rect 10704 7800 10732 7831
rect 10870 7828 10876 7880
rect 10928 7828 10934 7880
rect 11054 7828 11060 7880
rect 11112 7868 11118 7880
rect 11348 7877 11376 7976
rect 12342 7964 12348 7976
rect 12400 7964 12406 8016
rect 11606 7896 11612 7948
rect 11664 7896 11670 7948
rect 11333 7871 11391 7877
rect 11333 7868 11345 7871
rect 11112 7840 11345 7868
rect 11112 7828 11118 7840
rect 11333 7837 11345 7840
rect 11379 7837 11391 7871
rect 11333 7831 11391 7837
rect 11425 7871 11483 7877
rect 11425 7837 11437 7871
rect 11471 7868 11483 7871
rect 11624 7868 11652 7896
rect 11471 7840 11652 7868
rect 11471 7837 11483 7840
rect 11425 7831 11483 7837
rect 11440 7800 11468 7831
rect 11698 7828 11704 7880
rect 11756 7828 11762 7880
rect 10704 7772 11468 7800
rect 11609 7803 11667 7809
rect 9631 7769 9643 7772
rect 9585 7763 9643 7769
rect 11609 7769 11621 7803
rect 11655 7800 11667 7803
rect 11790 7800 11796 7812
rect 11655 7772 11796 7800
rect 11655 7769 11667 7772
rect 11609 7763 11667 7769
rect 11790 7760 11796 7772
rect 11848 7760 11854 7812
rect 4706 7692 4712 7744
rect 4764 7692 4770 7744
rect 5629 7735 5687 7741
rect 5629 7701 5641 7735
rect 5675 7732 5687 7735
rect 5902 7732 5908 7744
rect 5675 7704 5908 7732
rect 5675 7701 5687 7704
rect 5629 7695 5687 7701
rect 5902 7692 5908 7704
rect 5960 7692 5966 7744
rect 7282 7692 7288 7744
rect 7340 7732 7346 7744
rect 8297 7735 8355 7741
rect 8297 7732 8309 7735
rect 7340 7704 8309 7732
rect 7340 7692 7346 7704
rect 8297 7701 8309 7704
rect 8343 7701 8355 7735
rect 8297 7695 8355 7701
rect 8478 7692 8484 7744
rect 8536 7692 8542 7744
rect 9769 7735 9827 7741
rect 9769 7701 9781 7735
rect 9815 7732 9827 7735
rect 9858 7732 9864 7744
rect 9815 7704 9864 7732
rect 9815 7701 9827 7704
rect 9769 7695 9827 7701
rect 9858 7692 9864 7704
rect 9916 7692 9922 7744
rect 10778 7692 10784 7744
rect 10836 7732 10842 7744
rect 11054 7732 11060 7744
rect 10836 7704 11060 7732
rect 10836 7692 10842 7704
rect 11054 7692 11060 7704
rect 11112 7692 11118 7744
rect 11238 7692 11244 7744
rect 11296 7692 11302 7744
rect 11701 7735 11759 7741
rect 11701 7701 11713 7735
rect 11747 7732 11759 7735
rect 12250 7732 12256 7744
rect 11747 7704 12256 7732
rect 11747 7701 11759 7704
rect 11701 7695 11759 7701
rect 12250 7692 12256 7704
rect 12308 7692 12314 7744
rect 1104 7642 13708 7664
rect 1104 7590 3185 7642
rect 3237 7590 3249 7642
rect 3301 7590 3313 7642
rect 3365 7590 3377 7642
rect 3429 7590 3441 7642
rect 3493 7590 6336 7642
rect 6388 7590 6400 7642
rect 6452 7590 6464 7642
rect 6516 7590 6528 7642
rect 6580 7590 6592 7642
rect 6644 7590 9487 7642
rect 9539 7590 9551 7642
rect 9603 7590 9615 7642
rect 9667 7590 9679 7642
rect 9731 7590 9743 7642
rect 9795 7590 12638 7642
rect 12690 7590 12702 7642
rect 12754 7590 12766 7642
rect 12818 7590 12830 7642
rect 12882 7590 12894 7642
rect 12946 7590 13708 7642
rect 1104 7568 13708 7590
rect 4341 7531 4399 7537
rect 4341 7497 4353 7531
rect 4387 7528 4399 7531
rect 5166 7528 5172 7540
rect 4387 7500 5172 7528
rect 4387 7497 4399 7500
rect 4341 7491 4399 7497
rect 5166 7488 5172 7500
rect 5224 7488 5230 7540
rect 6457 7531 6515 7537
rect 6457 7528 6469 7531
rect 5736 7500 6469 7528
rect 2961 7463 3019 7469
rect 2961 7429 2973 7463
rect 3007 7460 3019 7463
rect 3007 7432 3648 7460
rect 3007 7429 3019 7432
rect 2961 7423 3019 7429
rect 3145 7395 3203 7401
rect 3145 7361 3157 7395
rect 3191 7392 3203 7395
rect 3191 7364 3372 7392
rect 3191 7361 3203 7364
rect 3145 7355 3203 7361
rect 2314 7148 2320 7200
rect 2372 7188 2378 7200
rect 3344 7197 3372 7364
rect 3510 7352 3516 7404
rect 3568 7352 3574 7404
rect 3620 7392 3648 7432
rect 3786 7420 3792 7472
rect 3844 7460 3850 7472
rect 4065 7463 4123 7469
rect 4065 7460 4077 7463
rect 3844 7432 4077 7460
rect 3844 7420 3850 7432
rect 4065 7429 4077 7432
rect 4111 7429 4123 7463
rect 5736 7460 5764 7500
rect 6457 7497 6469 7500
rect 6503 7497 6515 7531
rect 6457 7491 6515 7497
rect 6917 7531 6975 7537
rect 6917 7497 6929 7531
rect 6963 7528 6975 7531
rect 7190 7528 7196 7540
rect 6963 7500 7196 7528
rect 6963 7497 6975 7500
rect 6917 7491 6975 7497
rect 7190 7488 7196 7500
rect 7248 7488 7254 7540
rect 8570 7488 8576 7540
rect 8628 7528 8634 7540
rect 8846 7528 8852 7540
rect 8628 7500 8852 7528
rect 8628 7488 8634 7500
rect 8846 7488 8852 7500
rect 8904 7488 8910 7540
rect 9950 7528 9956 7540
rect 8956 7500 9956 7528
rect 5474 7432 5764 7460
rect 4065 7423 4123 7429
rect 5902 7420 5908 7472
rect 5960 7420 5966 7472
rect 6638 7460 6644 7472
rect 6564 7432 6644 7460
rect 3970 7392 3976 7404
rect 3620 7364 3976 7392
rect 3970 7352 3976 7364
rect 4028 7352 4034 7404
rect 6564 7401 6592 7432
rect 6638 7420 6644 7432
rect 6696 7460 6702 7472
rect 7098 7460 7104 7472
rect 6696 7432 7104 7460
rect 6696 7420 6702 7432
rect 7098 7420 7104 7432
rect 7156 7420 7162 7472
rect 8588 7460 8616 7488
rect 8665 7463 8723 7469
rect 8665 7460 8677 7463
rect 7300 7432 8677 7460
rect 4157 7395 4215 7401
rect 4157 7361 4169 7395
rect 4203 7392 4215 7395
rect 6549 7395 6607 7401
rect 4203 7364 4476 7392
rect 4203 7361 4215 7364
rect 4157 7355 4215 7361
rect 3697 7327 3755 7333
rect 3697 7293 3709 7327
rect 3743 7324 3755 7327
rect 3743 7296 3777 7324
rect 3743 7293 3755 7296
rect 3697 7287 3755 7293
rect 3602 7216 3608 7268
rect 3660 7256 3666 7268
rect 3712 7256 3740 7287
rect 3789 7259 3847 7265
rect 3789 7256 3801 7259
rect 3660 7228 3801 7256
rect 3660 7216 3666 7228
rect 3789 7225 3801 7228
rect 3835 7225 3847 7259
rect 3789 7219 3847 7225
rect 2777 7191 2835 7197
rect 2777 7188 2789 7191
rect 2372 7160 2789 7188
rect 2372 7148 2378 7160
rect 2777 7157 2789 7160
rect 2823 7157 2835 7191
rect 2777 7151 2835 7157
rect 3329 7191 3387 7197
rect 3329 7157 3341 7191
rect 3375 7188 3387 7191
rect 3694 7188 3700 7200
rect 3375 7160 3700 7188
rect 3375 7157 3387 7160
rect 3329 7151 3387 7157
rect 3694 7148 3700 7160
rect 3752 7148 3758 7200
rect 4448 7197 4476 7364
rect 6549 7361 6561 7395
rect 6595 7361 6607 7395
rect 6549 7355 6607 7361
rect 6730 7352 6736 7404
rect 6788 7392 6794 7404
rect 6825 7395 6883 7401
rect 6825 7392 6837 7395
rect 6788 7364 6837 7392
rect 6788 7352 6794 7364
rect 6825 7361 6837 7364
rect 6871 7392 6883 7395
rect 7300 7392 7328 7432
rect 8665 7429 8677 7432
rect 8711 7429 8723 7463
rect 8665 7423 8723 7429
rect 6871 7364 7328 7392
rect 6871 7361 6883 7364
rect 6825 7355 6883 7361
rect 7374 7352 7380 7404
rect 7432 7392 7438 7404
rect 8021 7395 8079 7401
rect 8021 7392 8033 7395
rect 7432 7364 8033 7392
rect 7432 7352 7438 7364
rect 8021 7361 8033 7364
rect 8067 7361 8079 7395
rect 8021 7355 8079 7361
rect 8570 7352 8576 7404
rect 8628 7392 8634 7404
rect 8956 7401 8984 7500
rect 9950 7488 9956 7500
rect 10008 7488 10014 7540
rect 11054 7488 11060 7540
rect 11112 7528 11118 7540
rect 11609 7531 11667 7537
rect 11609 7528 11621 7531
rect 11112 7500 11621 7528
rect 11112 7488 11118 7500
rect 11609 7497 11621 7500
rect 11655 7528 11667 7531
rect 11698 7528 11704 7540
rect 11655 7500 11704 7528
rect 11655 7497 11667 7500
rect 11609 7491 11667 7497
rect 11698 7488 11704 7500
rect 11756 7488 11762 7540
rect 11977 7531 12035 7537
rect 11977 7497 11989 7531
rect 12023 7528 12035 7531
rect 12269 7531 12327 7537
rect 12269 7528 12281 7531
rect 12023 7500 12281 7528
rect 12023 7497 12035 7500
rect 11977 7491 12035 7497
rect 12269 7497 12281 7500
rect 12315 7497 12327 7531
rect 12269 7491 12327 7497
rect 12437 7531 12495 7537
rect 12437 7497 12449 7531
rect 12483 7497 12495 7531
rect 12437 7491 12495 7497
rect 9769 7463 9827 7469
rect 9769 7429 9781 7463
rect 9815 7460 9827 7463
rect 9858 7460 9864 7472
rect 9815 7432 9864 7460
rect 9815 7429 9827 7432
rect 9769 7423 9827 7429
rect 9858 7420 9864 7432
rect 9916 7420 9922 7472
rect 11238 7460 11244 7472
rect 10994 7432 11244 7460
rect 11238 7420 11244 7432
rect 11296 7420 11302 7472
rect 12069 7463 12127 7469
rect 12069 7460 12081 7463
rect 11348 7432 12081 7460
rect 8849 7395 8907 7401
rect 8849 7392 8861 7395
rect 8628 7364 8861 7392
rect 8628 7352 8634 7364
rect 8849 7361 8861 7364
rect 8895 7361 8907 7395
rect 8849 7355 8907 7361
rect 8941 7395 8999 7401
rect 8941 7361 8953 7395
rect 8987 7361 8999 7395
rect 8941 7355 8999 7361
rect 9125 7395 9183 7401
rect 9125 7361 9137 7395
rect 9171 7392 9183 7395
rect 9398 7392 9404 7404
rect 9171 7364 9404 7392
rect 9171 7361 9183 7364
rect 9125 7355 9183 7361
rect 9398 7352 9404 7364
rect 9456 7352 9462 7404
rect 11348 7392 11376 7432
rect 12069 7429 12081 7432
rect 12115 7429 12127 7463
rect 12069 7423 12127 7429
rect 10980 7364 11376 7392
rect 6178 7284 6184 7336
rect 6236 7284 6242 7336
rect 8297 7327 8355 7333
rect 8297 7293 8309 7327
rect 8343 7293 8355 7327
rect 8297 7287 8355 7293
rect 8312 7256 8340 7287
rect 8662 7284 8668 7336
rect 8720 7324 8726 7336
rect 9033 7327 9091 7333
rect 9033 7324 9045 7327
rect 8720 7296 9045 7324
rect 8720 7284 8726 7296
rect 9033 7293 9045 7296
rect 9079 7293 9091 7327
rect 9033 7287 9091 7293
rect 9490 7284 9496 7336
rect 9548 7284 9554 7336
rect 10778 7324 10784 7336
rect 9600 7296 10784 7324
rect 9600 7256 9628 7296
rect 10778 7284 10784 7296
rect 10836 7284 10842 7336
rect 8312 7228 9628 7256
rect 4433 7191 4491 7197
rect 4433 7157 4445 7191
rect 4479 7188 4491 7191
rect 4614 7188 4620 7200
rect 4479 7160 4620 7188
rect 4479 7157 4491 7160
rect 4433 7151 4491 7157
rect 4614 7148 4620 7160
rect 4672 7148 4678 7200
rect 8846 7148 8852 7200
rect 8904 7188 8910 7200
rect 10502 7188 10508 7200
rect 8904 7160 10508 7188
rect 8904 7148 8910 7160
rect 10502 7148 10508 7160
rect 10560 7188 10566 7200
rect 10980 7188 11008 7364
rect 11422 7352 11428 7404
rect 11480 7392 11486 7404
rect 11517 7395 11575 7401
rect 11517 7392 11529 7395
rect 11480 7364 11529 7392
rect 11480 7352 11486 7364
rect 11517 7361 11529 7364
rect 11563 7392 11575 7395
rect 11606 7392 11612 7404
rect 11563 7364 11612 7392
rect 11563 7361 11575 7364
rect 11517 7355 11575 7361
rect 11606 7352 11612 7364
rect 11664 7352 11670 7404
rect 11790 7352 11796 7404
rect 11848 7352 11854 7404
rect 12452 7392 12480 7491
rect 12526 7420 12532 7472
rect 12584 7460 12590 7472
rect 12584 7432 13032 7460
rect 12584 7420 12590 7432
rect 13004 7401 13032 7432
rect 12713 7395 12771 7401
rect 12713 7392 12725 7395
rect 12452 7364 12725 7392
rect 12713 7361 12725 7364
rect 12759 7361 12771 7395
rect 12713 7355 12771 7361
rect 12989 7395 13047 7401
rect 12989 7361 13001 7395
rect 13035 7392 13047 7395
rect 13081 7395 13139 7401
rect 13081 7392 13093 7395
rect 13035 7364 13093 7392
rect 13035 7361 13047 7364
rect 12989 7355 13047 7361
rect 13081 7361 13093 7364
rect 13127 7361 13139 7395
rect 13081 7355 13139 7361
rect 11146 7284 11152 7336
rect 11204 7324 11210 7336
rect 11241 7327 11299 7333
rect 11241 7324 11253 7327
rect 11204 7296 11253 7324
rect 11204 7284 11210 7296
rect 11241 7293 11253 7296
rect 11287 7293 11299 7327
rect 11808 7324 11836 7352
rect 13262 7324 13268 7336
rect 11808 7296 13268 7324
rect 11241 7287 11299 7293
rect 13262 7284 13268 7296
rect 13320 7284 13326 7336
rect 10560 7160 11008 7188
rect 10560 7148 10566 7160
rect 12250 7148 12256 7200
rect 12308 7148 12314 7200
rect 12526 7148 12532 7200
rect 12584 7148 12590 7200
rect 12894 7148 12900 7200
rect 12952 7148 12958 7200
rect 13170 7148 13176 7200
rect 13228 7148 13234 7200
rect 1104 7098 13708 7120
rect 1104 7046 2525 7098
rect 2577 7046 2589 7098
rect 2641 7046 2653 7098
rect 2705 7046 2717 7098
rect 2769 7046 2781 7098
rect 2833 7046 5676 7098
rect 5728 7046 5740 7098
rect 5792 7046 5804 7098
rect 5856 7046 5868 7098
rect 5920 7046 5932 7098
rect 5984 7046 8827 7098
rect 8879 7046 8891 7098
rect 8943 7046 8955 7098
rect 9007 7046 9019 7098
rect 9071 7046 9083 7098
rect 9135 7046 11978 7098
rect 12030 7046 12042 7098
rect 12094 7046 12106 7098
rect 12158 7046 12170 7098
rect 12222 7046 12234 7098
rect 12286 7046 13708 7098
rect 1104 7024 13708 7046
rect 2314 6944 2320 6996
rect 2372 6944 2378 6996
rect 2777 6987 2835 6993
rect 2777 6953 2789 6987
rect 2823 6984 2835 6987
rect 2958 6984 2964 6996
rect 2823 6956 2964 6984
rect 2823 6953 2835 6956
rect 2777 6947 2835 6953
rect 2958 6944 2964 6956
rect 3016 6944 3022 6996
rect 4430 6984 4436 6996
rect 4080 6956 4436 6984
rect 2130 6876 2136 6928
rect 2188 6876 2194 6928
rect 2593 6919 2651 6925
rect 2593 6885 2605 6919
rect 2639 6885 2651 6919
rect 3326 6916 3332 6928
rect 2593 6879 2651 6885
rect 2746 6888 3332 6916
rect 2498 6848 2504 6860
rect 2056 6820 2504 6848
rect 1854 6740 1860 6792
rect 1912 6740 1918 6792
rect 2056 6789 2084 6820
rect 2498 6808 2504 6820
rect 2556 6808 2562 6860
rect 2041 6783 2099 6789
rect 2041 6749 2053 6783
rect 2087 6749 2099 6783
rect 2608 6780 2636 6879
rect 2746 6860 2774 6888
rect 3326 6876 3332 6888
rect 3384 6916 3390 6928
rect 3878 6916 3884 6928
rect 3384 6888 3884 6916
rect 3384 6876 3390 6888
rect 3878 6876 3884 6888
rect 3936 6876 3942 6928
rect 4080 6916 4108 6956
rect 4430 6944 4436 6956
rect 4488 6944 4494 6996
rect 7272 6987 7330 6993
rect 7272 6953 7284 6987
rect 7318 6984 7330 6987
rect 9306 6984 9312 6996
rect 7318 6956 9312 6984
rect 7318 6953 7330 6956
rect 7272 6947 7330 6953
rect 9306 6944 9312 6956
rect 9364 6944 9370 6996
rect 9674 6944 9680 6996
rect 9732 6984 9738 6996
rect 10318 6984 10324 6996
rect 9732 6956 10324 6984
rect 9732 6944 9738 6956
rect 10318 6944 10324 6956
rect 10376 6944 10382 6996
rect 10413 6987 10471 6993
rect 10413 6953 10425 6987
rect 10459 6984 10471 6987
rect 11238 6984 11244 6996
rect 10459 6956 11244 6984
rect 10459 6953 10471 6956
rect 10413 6947 10471 6953
rect 11238 6944 11244 6956
rect 11296 6944 11302 6996
rect 11780 6987 11838 6993
rect 11780 6953 11792 6987
rect 11826 6984 11838 6987
rect 12526 6984 12532 6996
rect 11826 6956 12532 6984
rect 11826 6953 11838 6956
rect 11780 6947 11838 6953
rect 12526 6944 12532 6956
rect 12584 6944 12590 6996
rect 3988 6888 4108 6916
rect 2682 6808 2688 6860
rect 2740 6820 2774 6860
rect 3237 6851 3295 6857
rect 2740 6808 2746 6820
rect 3237 6817 3249 6851
rect 3283 6848 3295 6851
rect 3602 6848 3608 6860
rect 3283 6820 3608 6848
rect 3283 6817 3295 6820
rect 3237 6811 3295 6817
rect 3602 6808 3608 6820
rect 3660 6808 3666 6860
rect 3988 6848 4016 6888
rect 8294 6876 8300 6928
rect 8352 6916 8358 6928
rect 8846 6916 8852 6928
rect 8352 6888 8852 6916
rect 8352 6876 8358 6888
rect 8846 6876 8852 6888
rect 8904 6876 8910 6928
rect 9214 6876 9220 6928
rect 9272 6916 9278 6928
rect 10686 6916 10692 6928
rect 9272 6888 10692 6916
rect 9272 6876 9278 6888
rect 10686 6876 10692 6888
rect 10744 6876 10750 6928
rect 3712 6820 4016 6848
rect 2041 6743 2099 6749
rect 2424 6752 2636 6780
rect 3145 6783 3203 6789
rect 1486 6672 1492 6724
rect 1544 6712 1550 6724
rect 2424 6712 2452 6752
rect 3145 6749 3157 6783
rect 3191 6749 3203 6783
rect 3145 6743 3203 6749
rect 1544 6684 2452 6712
rect 2501 6715 2559 6721
rect 1544 6672 1550 6684
rect 2501 6681 2513 6715
rect 2547 6712 2559 6715
rect 2961 6715 3019 6721
rect 2961 6712 2973 6715
rect 2547 6684 2973 6712
rect 2547 6681 2559 6684
rect 2501 6675 2559 6681
rect 2961 6681 2973 6684
rect 3007 6712 3019 6715
rect 3050 6712 3056 6724
rect 3007 6684 3056 6712
rect 3007 6681 3019 6684
rect 2961 6675 3019 6681
rect 3050 6672 3056 6684
rect 3108 6672 3114 6724
rect 3160 6712 3188 6743
rect 3326 6740 3332 6792
rect 3384 6740 3390 6792
rect 3421 6783 3479 6789
rect 3421 6749 3433 6783
rect 3467 6780 3479 6783
rect 3510 6780 3516 6792
rect 3467 6752 3516 6780
rect 3467 6749 3479 6752
rect 3421 6743 3479 6749
rect 3510 6740 3516 6752
rect 3568 6780 3574 6792
rect 3712 6780 3740 6820
rect 4062 6808 4068 6860
rect 4120 6848 4126 6860
rect 4890 6848 4896 6860
rect 4120 6820 4896 6848
rect 4120 6808 4126 6820
rect 4890 6808 4896 6820
rect 4948 6808 4954 6860
rect 6638 6808 6644 6860
rect 6696 6808 6702 6860
rect 7009 6851 7067 6857
rect 7009 6817 7021 6851
rect 7055 6848 7067 6851
rect 9490 6848 9496 6860
rect 7055 6820 9496 6848
rect 7055 6817 7067 6820
rect 7009 6811 7067 6817
rect 9490 6808 9496 6820
rect 9548 6848 9554 6860
rect 10410 6848 10416 6860
rect 9548 6820 10416 6848
rect 9548 6808 9554 6820
rect 10410 6808 10416 6820
rect 10468 6848 10474 6860
rect 11517 6851 11575 6857
rect 11517 6848 11529 6851
rect 10468 6820 11529 6848
rect 10468 6808 10474 6820
rect 11517 6817 11529 6820
rect 11563 6817 11575 6851
rect 11517 6811 11575 6817
rect 13262 6808 13268 6860
rect 13320 6808 13326 6860
rect 3568 6752 3740 6780
rect 3568 6740 3574 6752
rect 3786 6740 3792 6792
rect 3844 6740 3850 6792
rect 3970 6740 3976 6792
rect 4028 6740 4034 6792
rect 6089 6783 6147 6789
rect 6089 6749 6101 6783
rect 6135 6780 6147 6783
rect 6656 6780 6684 6808
rect 6135 6752 6684 6780
rect 6917 6783 6975 6789
rect 6135 6749 6147 6752
rect 6089 6743 6147 6749
rect 6917 6749 6929 6783
rect 6963 6749 6975 6783
rect 6917 6743 6975 6749
rect 3804 6712 3832 6740
rect 3160 6684 4292 6712
rect 2041 6647 2099 6653
rect 2041 6613 2053 6647
rect 2087 6644 2099 6647
rect 2291 6647 2349 6653
rect 2291 6644 2303 6647
rect 2087 6616 2303 6644
rect 2087 6613 2099 6616
rect 2041 6607 2099 6613
rect 2291 6613 2303 6616
rect 2337 6613 2349 6647
rect 2291 6607 2349 6613
rect 2761 6647 2819 6653
rect 2761 6613 2773 6647
rect 2807 6644 2819 6647
rect 3510 6644 3516 6656
rect 2807 6616 3516 6644
rect 2807 6613 2819 6616
rect 2761 6607 2819 6613
rect 3510 6604 3516 6616
rect 3568 6604 3574 6656
rect 3605 6647 3663 6653
rect 3605 6613 3617 6647
rect 3651 6644 3663 6647
rect 3878 6644 3884 6656
rect 3651 6616 3884 6644
rect 3651 6613 3663 6616
rect 3605 6607 3663 6613
rect 3878 6604 3884 6616
rect 3936 6604 3942 6656
rect 3973 6647 4031 6653
rect 3973 6613 3985 6647
rect 4019 6644 4031 6647
rect 4154 6644 4160 6656
rect 4019 6616 4160 6644
rect 4019 6613 4031 6616
rect 3973 6607 4031 6613
rect 4154 6604 4160 6616
rect 4212 6604 4218 6656
rect 4264 6644 4292 6684
rect 4338 6672 4344 6724
rect 4396 6672 4402 6724
rect 5997 6715 6055 6721
rect 5997 6712 6009 6715
rect 5566 6684 6009 6712
rect 5997 6681 6009 6684
rect 6043 6681 6055 6715
rect 6932 6712 6960 6743
rect 9214 6740 9220 6792
rect 9272 6740 9278 6792
rect 10042 6740 10048 6792
rect 10100 6740 10106 6792
rect 10134 6740 10140 6792
rect 10192 6740 10198 6792
rect 10226 6740 10232 6792
rect 10284 6780 10290 6792
rect 10778 6780 10784 6792
rect 10284 6752 10784 6780
rect 10284 6740 10290 6752
rect 10778 6740 10784 6752
rect 10836 6740 10842 6792
rect 10870 6740 10876 6792
rect 10928 6740 10934 6792
rect 11241 6783 11299 6789
rect 11241 6780 11253 6783
rect 10980 6752 11253 6780
rect 7374 6712 7380 6724
rect 6932 6684 7380 6712
rect 5997 6675 6055 6681
rect 7374 6672 7380 6684
rect 7432 6672 7438 6724
rect 8294 6672 8300 6724
rect 8352 6672 8358 6724
rect 9232 6712 9260 6740
rect 8772 6684 9260 6712
rect 9769 6715 9827 6721
rect 5810 6644 5816 6656
rect 4264 6616 5816 6644
rect 5810 6604 5816 6616
rect 5868 6604 5874 6656
rect 8772 6653 8800 6684
rect 9769 6681 9781 6715
rect 9815 6712 9827 6715
rect 10505 6715 10563 6721
rect 9815 6684 10088 6712
rect 9815 6681 9827 6684
rect 9769 6675 9827 6681
rect 10060 6656 10088 6684
rect 10505 6681 10517 6715
rect 10551 6712 10563 6715
rect 10980 6712 11008 6752
rect 11241 6749 11253 6752
rect 11287 6780 11299 6783
rect 11422 6780 11428 6792
rect 11287 6752 11428 6780
rect 11287 6749 11299 6752
rect 11241 6743 11299 6749
rect 11422 6740 11428 6752
rect 11480 6740 11486 6792
rect 12894 6740 12900 6792
rect 12952 6740 12958 6792
rect 10551 6684 11008 6712
rect 11149 6715 11207 6721
rect 10551 6681 10563 6684
rect 10505 6675 10563 6681
rect 11149 6681 11161 6715
rect 11195 6712 11207 6715
rect 11330 6712 11336 6724
rect 11195 6684 11336 6712
rect 11195 6681 11207 6684
rect 11149 6675 11207 6681
rect 11330 6672 11336 6684
rect 11388 6672 11394 6724
rect 8757 6647 8815 6653
rect 8757 6613 8769 6647
rect 8803 6613 8815 6647
rect 8757 6607 8815 6613
rect 9030 6604 9036 6656
rect 9088 6644 9094 6656
rect 9674 6644 9680 6656
rect 9088 6616 9680 6644
rect 9088 6604 9094 6616
rect 9674 6604 9680 6616
rect 9732 6604 9738 6656
rect 9858 6604 9864 6656
rect 9916 6604 9922 6656
rect 10042 6604 10048 6656
rect 10100 6604 10106 6656
rect 10594 6604 10600 6656
rect 10652 6604 10658 6656
rect 11054 6604 11060 6656
rect 11112 6604 11118 6656
rect 1104 6554 13708 6576
rect 1104 6502 3185 6554
rect 3237 6502 3249 6554
rect 3301 6502 3313 6554
rect 3365 6502 3377 6554
rect 3429 6502 3441 6554
rect 3493 6502 6336 6554
rect 6388 6502 6400 6554
rect 6452 6502 6464 6554
rect 6516 6502 6528 6554
rect 6580 6502 6592 6554
rect 6644 6502 9487 6554
rect 9539 6502 9551 6554
rect 9603 6502 9615 6554
rect 9667 6502 9679 6554
rect 9731 6502 9743 6554
rect 9795 6502 12638 6554
rect 12690 6502 12702 6554
rect 12754 6502 12766 6554
rect 12818 6502 12830 6554
rect 12882 6502 12894 6554
rect 12946 6502 13708 6554
rect 1104 6480 13708 6502
rect 4062 6440 4068 6452
rect 1872 6412 4068 6440
rect 1872 6372 1900 6412
rect 4062 6400 4068 6412
rect 4120 6400 4126 6452
rect 4338 6400 4344 6452
rect 4396 6440 4402 6452
rect 4433 6443 4491 6449
rect 4433 6440 4445 6443
rect 4396 6412 4445 6440
rect 4396 6400 4402 6412
rect 4433 6409 4445 6412
rect 4479 6409 4491 6443
rect 4433 6403 4491 6409
rect 4706 6400 4712 6452
rect 4764 6440 4770 6452
rect 5077 6443 5135 6449
rect 5077 6440 5089 6443
rect 4764 6412 5089 6440
rect 4764 6400 4770 6412
rect 5077 6409 5089 6412
rect 5123 6409 5135 6443
rect 5077 6403 5135 6409
rect 6641 6443 6699 6449
rect 6641 6409 6653 6443
rect 6687 6409 6699 6443
rect 6641 6403 6699 6409
rect 8205 6443 8263 6449
rect 8205 6409 8217 6443
rect 8251 6440 8263 6443
rect 8294 6440 8300 6452
rect 8251 6412 8300 6440
rect 8251 6409 8263 6412
rect 8205 6403 8263 6409
rect 1780 6344 1900 6372
rect 1780 6316 1808 6344
rect 3050 6332 3056 6384
rect 3108 6332 3114 6384
rect 4522 6372 4528 6384
rect 3804 6344 4528 6372
rect 1486 6264 1492 6316
rect 1544 6264 1550 6316
rect 1762 6264 1768 6316
rect 1820 6264 1826 6316
rect 3804 6313 3832 6344
rect 4522 6332 4528 6344
rect 4580 6372 4586 6384
rect 6086 6372 6092 6384
rect 4580 6344 6092 6372
rect 4580 6332 4586 6344
rect 6086 6332 6092 6344
rect 6144 6372 6150 6384
rect 6656 6372 6684 6403
rect 8294 6400 8300 6412
rect 8352 6400 8358 6452
rect 9030 6400 9036 6452
rect 9088 6440 9094 6452
rect 9088 6412 9260 6440
rect 9088 6400 9094 6412
rect 9048 6372 9076 6400
rect 6144 6344 9076 6372
rect 6144 6332 6150 6344
rect 3789 6307 3847 6313
rect 3789 6273 3801 6307
rect 3835 6273 3847 6307
rect 3789 6267 3847 6273
rect 3878 6264 3884 6316
rect 3936 6304 3942 6316
rect 3973 6307 4031 6313
rect 3973 6304 3985 6307
rect 3936 6276 3985 6304
rect 3936 6264 3942 6276
rect 3973 6273 3985 6276
rect 4019 6273 4031 6307
rect 3973 6267 4031 6273
rect 4065 6307 4123 6313
rect 4065 6273 4077 6307
rect 4111 6273 4123 6307
rect 4065 6267 4123 6273
rect 2041 6239 2099 6245
rect 2041 6236 2053 6239
rect 1688 6208 2053 6236
rect 1688 6177 1716 6208
rect 2041 6205 2053 6208
rect 2087 6205 2099 6239
rect 2041 6199 2099 6205
rect 3418 6196 3424 6248
rect 3476 6236 3482 6248
rect 4080 6236 4108 6267
rect 4154 6264 4160 6316
rect 4212 6264 4218 6316
rect 4614 6264 4620 6316
rect 4672 6264 4678 6316
rect 4801 6307 4859 6313
rect 4801 6273 4813 6307
rect 4847 6304 4859 6307
rect 5810 6304 5816 6316
rect 4847 6276 5816 6304
rect 4847 6273 4859 6276
rect 4801 6267 4859 6273
rect 5810 6264 5816 6276
rect 5868 6264 5874 6316
rect 6457 6307 6515 6313
rect 6457 6273 6469 6307
rect 6503 6304 6515 6307
rect 6730 6304 6736 6316
rect 6503 6276 6736 6304
rect 6503 6273 6515 6276
rect 6457 6267 6515 6273
rect 6730 6264 6736 6276
rect 6788 6264 6794 6316
rect 7374 6264 7380 6316
rect 7432 6304 7438 6316
rect 8021 6307 8079 6313
rect 8021 6304 8033 6307
rect 7432 6276 8033 6304
rect 7432 6264 7438 6276
rect 8021 6273 8033 6276
rect 8067 6304 8079 6307
rect 8113 6307 8171 6313
rect 8113 6304 8125 6307
rect 8067 6276 8125 6304
rect 8067 6273 8079 6276
rect 8021 6267 8079 6273
rect 8113 6273 8125 6276
rect 8159 6273 8171 6307
rect 8113 6267 8171 6273
rect 8665 6307 8723 6313
rect 8665 6273 8677 6307
rect 8711 6304 8723 6307
rect 8846 6304 8852 6316
rect 8711 6276 8852 6304
rect 8711 6273 8723 6276
rect 8665 6267 8723 6273
rect 8846 6264 8852 6276
rect 8904 6264 8910 6316
rect 9232 6313 9260 6412
rect 9306 6400 9312 6452
rect 9364 6440 9370 6452
rect 9493 6443 9551 6449
rect 9493 6440 9505 6443
rect 9364 6412 9505 6440
rect 9364 6400 9370 6412
rect 9493 6409 9505 6412
rect 9539 6409 9551 6443
rect 9769 6443 9827 6449
rect 9769 6440 9781 6443
rect 9493 6403 9551 6409
rect 9600 6412 9781 6440
rect 9398 6332 9404 6384
rect 9456 6372 9462 6384
rect 9600 6372 9628 6412
rect 9769 6409 9781 6412
rect 9815 6409 9827 6443
rect 9769 6403 9827 6409
rect 9858 6400 9864 6452
rect 9916 6440 9922 6452
rect 10613 6443 10671 6449
rect 10613 6440 10625 6443
rect 9916 6412 10625 6440
rect 9916 6400 9922 6412
rect 10613 6409 10625 6412
rect 10659 6409 10671 6443
rect 10613 6403 10671 6409
rect 11238 6400 11244 6452
rect 11296 6400 11302 6452
rect 13265 6443 13323 6449
rect 13265 6440 13277 6443
rect 11348 6412 13277 6440
rect 10226 6372 10232 6384
rect 9456 6344 9628 6372
rect 9968 6344 10232 6372
rect 9456 6332 9462 6344
rect 9125 6307 9183 6313
rect 9125 6273 9137 6307
rect 9171 6273 9183 6307
rect 9125 6267 9183 6273
rect 9217 6307 9275 6313
rect 9217 6273 9229 6307
rect 9263 6273 9275 6307
rect 9217 6267 9275 6273
rect 3476 6208 4108 6236
rect 3476 6196 3482 6208
rect 4246 6196 4252 6248
rect 4304 6236 4310 6248
rect 4709 6239 4767 6245
rect 4709 6236 4721 6239
rect 4304 6208 4721 6236
rect 4304 6196 4310 6208
rect 4709 6205 4721 6208
rect 4755 6205 4767 6239
rect 4709 6199 4767 6205
rect 4893 6239 4951 6245
rect 4893 6205 4905 6239
rect 4939 6205 4951 6239
rect 4893 6199 4951 6205
rect 7837 6239 7895 6245
rect 7837 6205 7849 6239
rect 7883 6236 7895 6239
rect 7926 6236 7932 6248
rect 7883 6208 7932 6236
rect 7883 6205 7895 6208
rect 7837 6199 7895 6205
rect 1673 6171 1731 6177
rect 1673 6137 1685 6171
rect 1719 6137 1731 6171
rect 3694 6168 3700 6180
rect 1673 6131 1731 6137
rect 3436 6140 3700 6168
rect 1854 6060 1860 6112
rect 1912 6100 1918 6112
rect 3436 6100 3464 6140
rect 3694 6128 3700 6140
rect 3752 6168 3758 6180
rect 4908 6168 4936 6199
rect 7926 6196 7932 6208
rect 7984 6196 7990 6248
rect 8386 6196 8392 6248
rect 8444 6236 8450 6248
rect 8757 6239 8815 6245
rect 8757 6236 8769 6239
rect 8444 6208 8769 6236
rect 8444 6196 8450 6208
rect 8757 6205 8769 6208
rect 8803 6205 8815 6239
rect 9140 6236 9168 6267
rect 9582 6264 9588 6316
rect 9640 6264 9646 6316
rect 9674 6264 9680 6316
rect 9732 6264 9738 6316
rect 9968 6313 9996 6344
rect 10226 6332 10232 6344
rect 10284 6332 10290 6384
rect 10413 6375 10471 6381
rect 10413 6341 10425 6375
rect 10459 6372 10471 6375
rect 10502 6372 10508 6384
rect 10459 6344 10508 6372
rect 10459 6341 10471 6344
rect 10413 6335 10471 6341
rect 10502 6332 10508 6344
rect 10560 6332 10566 6384
rect 10778 6332 10784 6384
rect 10836 6372 10842 6384
rect 11348 6372 11376 6412
rect 13265 6409 13277 6412
rect 13311 6409 13323 6443
rect 13265 6403 13323 6409
rect 13170 6372 13176 6384
rect 10836 6344 11376 6372
rect 13018 6344 13176 6372
rect 10836 6332 10842 6344
rect 9777 6305 9835 6311
rect 9777 6271 9789 6305
rect 9823 6302 9835 6305
rect 9953 6307 10011 6313
rect 9823 6274 9904 6302
rect 9823 6271 9835 6274
rect 9777 6265 9835 6271
rect 9677 6259 9689 6264
rect 9723 6259 9735 6264
rect 9677 6253 9735 6259
rect 9306 6236 9312 6248
rect 9140 6208 9312 6236
rect 8757 6199 8815 6205
rect 9306 6196 9312 6208
rect 9364 6196 9370 6248
rect 9876 6236 9904 6274
rect 9953 6273 9965 6307
rect 9999 6273 10011 6307
rect 9953 6267 10011 6273
rect 10042 6264 10048 6316
rect 10100 6264 10106 6316
rect 10686 6304 10692 6316
rect 10152 6276 10692 6304
rect 10152 6236 10180 6276
rect 10686 6264 10692 6276
rect 10744 6304 10750 6316
rect 10873 6307 10931 6313
rect 10873 6304 10885 6307
rect 10744 6276 10885 6304
rect 10744 6264 10750 6276
rect 10873 6273 10885 6276
rect 10919 6273 10931 6307
rect 10873 6267 10931 6273
rect 11054 6264 11060 6316
rect 11112 6264 11118 6316
rect 11348 6313 11376 6344
rect 13170 6332 13176 6344
rect 13228 6332 13234 6384
rect 11333 6307 11391 6313
rect 11333 6273 11345 6307
rect 11379 6273 11391 6307
rect 11333 6267 11391 6273
rect 9876 6208 10180 6236
rect 10502 6196 10508 6248
rect 10560 6236 10566 6248
rect 11517 6239 11575 6245
rect 11517 6236 11529 6239
rect 10560 6208 11529 6236
rect 10560 6196 10566 6208
rect 11517 6205 11529 6208
rect 11563 6205 11575 6239
rect 11517 6199 11575 6205
rect 11790 6196 11796 6248
rect 11848 6196 11854 6248
rect 3752 6140 4936 6168
rect 3752 6128 3758 6140
rect 8662 6128 8668 6180
rect 8720 6168 8726 6180
rect 10965 6171 11023 6177
rect 10965 6168 10977 6171
rect 8720 6140 10977 6168
rect 8720 6128 8726 6140
rect 1912 6072 3464 6100
rect 3513 6103 3571 6109
rect 1912 6060 1918 6072
rect 3513 6069 3525 6103
rect 3559 6100 3571 6103
rect 3602 6100 3608 6112
rect 3559 6072 3608 6100
rect 3559 6069 3571 6072
rect 3513 6063 3571 6069
rect 3602 6060 3608 6072
rect 3660 6100 3666 6112
rect 3970 6100 3976 6112
rect 3660 6072 3976 6100
rect 3660 6060 3666 6072
rect 3970 6060 3976 6072
rect 4028 6060 4034 6112
rect 8478 6060 8484 6112
rect 8536 6060 8542 6112
rect 9048 6109 9076 6140
rect 10965 6137 10977 6140
rect 11011 6137 11023 6171
rect 10965 6131 11023 6137
rect 9033 6103 9091 6109
rect 9033 6069 9045 6103
rect 9079 6069 9091 6103
rect 9033 6063 9091 6069
rect 9582 6060 9588 6112
rect 9640 6100 9646 6112
rect 10137 6103 10195 6109
rect 10137 6100 10149 6103
rect 9640 6072 10149 6100
rect 9640 6060 9646 6072
rect 10137 6069 10149 6072
rect 10183 6069 10195 6103
rect 10137 6063 10195 6069
rect 10594 6060 10600 6112
rect 10652 6060 10658 6112
rect 10778 6060 10784 6112
rect 10836 6060 10842 6112
rect 1104 6010 13708 6032
rect 1104 5958 2525 6010
rect 2577 5958 2589 6010
rect 2641 5958 2653 6010
rect 2705 5958 2717 6010
rect 2769 5958 2781 6010
rect 2833 5958 5676 6010
rect 5728 5958 5740 6010
rect 5792 5958 5804 6010
rect 5856 5958 5868 6010
rect 5920 5958 5932 6010
rect 5984 5958 8827 6010
rect 8879 5958 8891 6010
rect 8943 5958 8955 6010
rect 9007 5958 9019 6010
rect 9071 5958 9083 6010
rect 9135 5958 11978 6010
rect 12030 5958 12042 6010
rect 12094 5958 12106 6010
rect 12158 5958 12170 6010
rect 12222 5958 12234 6010
rect 12286 5958 13708 6010
rect 1104 5936 13708 5958
rect 3510 5856 3516 5908
rect 3568 5896 3574 5908
rect 3789 5899 3847 5905
rect 3789 5896 3801 5899
rect 3568 5868 3801 5896
rect 3568 5856 3574 5868
rect 3789 5865 3801 5868
rect 3835 5865 3847 5899
rect 3789 5859 3847 5865
rect 4890 5856 4896 5908
rect 4948 5896 4954 5908
rect 5261 5899 5319 5905
rect 5261 5896 5273 5899
rect 4948 5868 5273 5896
rect 4948 5856 4954 5868
rect 5261 5865 5273 5868
rect 5307 5896 5319 5899
rect 6178 5896 6184 5908
rect 5307 5868 6184 5896
rect 5307 5865 5319 5868
rect 5261 5859 5319 5865
rect 6178 5856 6184 5868
rect 6236 5856 6242 5908
rect 10410 5856 10416 5908
rect 10468 5856 10474 5908
rect 11333 5899 11391 5905
rect 11333 5865 11345 5899
rect 11379 5896 11391 5899
rect 11790 5896 11796 5908
rect 11379 5868 11796 5896
rect 11379 5865 11391 5868
rect 11333 5859 11391 5865
rect 11790 5856 11796 5868
rect 11848 5856 11854 5908
rect 3237 5831 3295 5837
rect 3237 5797 3249 5831
rect 3283 5828 3295 5831
rect 4062 5828 4068 5840
rect 3283 5800 4068 5828
rect 3283 5797 3295 5800
rect 3237 5791 3295 5797
rect 4062 5788 4068 5800
rect 4120 5788 4126 5840
rect 1489 5763 1547 5769
rect 1489 5729 1501 5763
rect 1535 5760 1547 5763
rect 1762 5760 1768 5772
rect 1535 5732 1768 5760
rect 1535 5729 1547 5732
rect 1489 5723 1547 5729
rect 1762 5720 1768 5732
rect 1820 5720 1826 5772
rect 2958 5720 2964 5772
rect 3016 5760 3022 5772
rect 3418 5760 3424 5772
rect 3016 5732 3424 5760
rect 3016 5720 3022 5732
rect 3418 5720 3424 5732
rect 3476 5760 3482 5772
rect 3513 5763 3571 5769
rect 3513 5760 3525 5763
rect 3476 5732 3525 5760
rect 3476 5720 3482 5732
rect 3513 5729 3525 5732
rect 3559 5729 3571 5763
rect 3513 5723 3571 5729
rect 2866 5652 2872 5704
rect 2924 5652 2930 5704
rect 3605 5695 3663 5701
rect 3605 5661 3617 5695
rect 3651 5692 3663 5695
rect 3694 5692 3700 5704
rect 3651 5664 3700 5692
rect 3651 5661 3663 5664
rect 3605 5655 3663 5661
rect 3694 5652 3700 5664
rect 3752 5652 3758 5704
rect 3970 5652 3976 5704
rect 4028 5652 4034 5704
rect 6549 5695 6607 5701
rect 6549 5661 6561 5695
rect 6595 5692 6607 5695
rect 6822 5692 6828 5704
rect 6595 5664 6828 5692
rect 6595 5661 6607 5664
rect 6549 5655 6607 5661
rect 6822 5652 6828 5664
rect 6880 5692 6886 5704
rect 9125 5695 9183 5701
rect 9125 5692 9137 5695
rect 6880 5664 9137 5692
rect 6880 5652 6886 5664
rect 9125 5661 9137 5664
rect 9171 5661 9183 5695
rect 9125 5655 9183 5661
rect 10778 5652 10784 5704
rect 10836 5692 10842 5704
rect 11149 5695 11207 5701
rect 11149 5692 11161 5695
rect 10836 5664 11161 5692
rect 10836 5652 10842 5664
rect 11149 5661 11161 5664
rect 11195 5661 11207 5695
rect 11149 5655 11207 5661
rect 1762 5584 1768 5636
rect 1820 5584 1826 5636
rect 4157 5627 4215 5633
rect 4157 5593 4169 5627
rect 4203 5624 4215 5627
rect 4246 5624 4252 5636
rect 4203 5596 4252 5624
rect 4203 5593 4215 5596
rect 4157 5587 4215 5593
rect 4246 5584 4252 5596
rect 4304 5584 4310 5636
rect 1104 5466 13708 5488
rect 1104 5414 3185 5466
rect 3237 5414 3249 5466
rect 3301 5414 3313 5466
rect 3365 5414 3377 5466
rect 3429 5414 3441 5466
rect 3493 5414 6336 5466
rect 6388 5414 6400 5466
rect 6452 5414 6464 5466
rect 6516 5414 6528 5466
rect 6580 5414 6592 5466
rect 6644 5414 9487 5466
rect 9539 5414 9551 5466
rect 9603 5414 9615 5466
rect 9667 5414 9679 5466
rect 9731 5414 9743 5466
rect 9795 5414 12638 5466
rect 12690 5414 12702 5466
rect 12754 5414 12766 5466
rect 12818 5414 12830 5466
rect 12882 5414 12894 5466
rect 12946 5414 13708 5466
rect 1104 5392 13708 5414
rect 1762 5312 1768 5364
rect 1820 5352 1826 5364
rect 2133 5355 2191 5361
rect 2133 5352 2145 5355
rect 1820 5324 2145 5352
rect 1820 5312 1826 5324
rect 2133 5321 2145 5324
rect 2179 5321 2191 5355
rect 2133 5315 2191 5321
rect 2961 5355 3019 5361
rect 2961 5321 2973 5355
rect 3007 5352 3019 5355
rect 3050 5352 3056 5364
rect 3007 5324 3056 5352
rect 3007 5321 3019 5324
rect 2961 5315 3019 5321
rect 3050 5312 3056 5324
rect 3108 5312 3114 5364
rect 2866 5244 2872 5296
rect 2924 5284 2930 5296
rect 3237 5287 3295 5293
rect 3237 5284 3249 5287
rect 2924 5256 3249 5284
rect 2924 5244 2930 5256
rect 3237 5253 3249 5256
rect 3283 5253 3295 5287
rect 3237 5247 3295 5253
rect 4890 5244 4896 5296
rect 4948 5244 4954 5296
rect 2130 5176 2136 5228
rect 2188 5216 2194 5228
rect 2317 5219 2375 5225
rect 2317 5216 2329 5219
rect 2188 5188 2329 5216
rect 2188 5176 2194 5188
rect 2317 5185 2329 5188
rect 2363 5185 2375 5219
rect 2317 5179 2375 5185
rect 3053 5219 3111 5225
rect 3053 5185 3065 5219
rect 3099 5216 3111 5219
rect 3329 5219 3387 5225
rect 3329 5216 3341 5219
rect 3099 5188 3341 5216
rect 3099 5185 3111 5188
rect 3053 5179 3111 5185
rect 3329 5185 3341 5188
rect 3375 5216 3387 5219
rect 3602 5216 3608 5228
rect 3375 5188 3608 5216
rect 3375 5185 3387 5188
rect 3329 5179 3387 5185
rect 3602 5176 3608 5188
rect 3660 5176 3666 5228
rect 5534 5108 5540 5160
rect 5592 5108 5598 5160
rect 5905 5083 5963 5089
rect 5905 5049 5917 5083
rect 5951 5080 5963 5083
rect 6086 5080 6092 5092
rect 5951 5052 6092 5080
rect 5951 5049 5963 5052
rect 5905 5043 5963 5049
rect 6086 5040 6092 5052
rect 6144 5040 6150 5092
rect 5994 4972 6000 5024
rect 6052 4972 6058 5024
rect 9674 4972 9680 5024
rect 9732 5012 9738 5024
rect 10778 5012 10784 5024
rect 9732 4984 10784 5012
rect 9732 4972 9738 4984
rect 10778 4972 10784 4984
rect 10836 4972 10842 5024
rect 1104 4922 13708 4944
rect 1104 4870 2525 4922
rect 2577 4870 2589 4922
rect 2641 4870 2653 4922
rect 2705 4870 2717 4922
rect 2769 4870 2781 4922
rect 2833 4870 5676 4922
rect 5728 4870 5740 4922
rect 5792 4870 5804 4922
rect 5856 4870 5868 4922
rect 5920 4870 5932 4922
rect 5984 4870 8827 4922
rect 8879 4870 8891 4922
rect 8943 4870 8955 4922
rect 9007 4870 9019 4922
rect 9071 4870 9083 4922
rect 9135 4870 11978 4922
rect 12030 4870 12042 4922
rect 12094 4870 12106 4922
rect 12158 4870 12170 4922
rect 12222 4870 12234 4922
rect 12286 4870 13708 4922
rect 1104 4848 13708 4870
rect 3970 4768 3976 4820
rect 4028 4808 4034 4820
rect 4798 4808 4804 4820
rect 4028 4780 4804 4808
rect 4028 4768 4034 4780
rect 4798 4768 4804 4780
rect 4856 4768 4862 4820
rect 7926 4808 7932 4820
rect 4908 4780 7932 4808
rect 3602 4700 3608 4752
rect 3660 4740 3666 4752
rect 4908 4740 4936 4780
rect 3660 4712 4936 4740
rect 3660 4700 3666 4712
rect 6822 4700 6828 4752
rect 6880 4740 6886 4752
rect 7193 4743 7251 4749
rect 7193 4740 7205 4743
rect 6880 4712 7205 4740
rect 6880 4700 6886 4712
rect 7193 4709 7205 4712
rect 7239 4709 7251 4743
rect 7193 4703 7251 4709
rect 4062 4632 4068 4684
rect 4120 4672 4126 4684
rect 4890 4672 4896 4684
rect 4120 4644 4896 4672
rect 4120 4632 4126 4644
rect 4890 4632 4896 4644
rect 4948 4672 4954 4684
rect 5442 4672 5448 4684
rect 4948 4644 5448 4672
rect 4948 4632 4954 4644
rect 5442 4632 5448 4644
rect 5500 4632 5506 4684
rect 4338 4564 4344 4616
rect 4396 4564 4402 4616
rect 4798 4564 4804 4616
rect 4856 4604 4862 4616
rect 7484 4613 7512 4780
rect 7926 4768 7932 4780
rect 7984 4808 7990 4820
rect 7984 4780 12434 4808
rect 7984 4768 7990 4780
rect 9416 4712 10456 4740
rect 8570 4672 8576 4684
rect 8404 4644 8576 4672
rect 8404 4613 8432 4644
rect 8570 4632 8576 4644
rect 8628 4672 8634 4684
rect 9416 4681 9444 4712
rect 9401 4675 9459 4681
rect 9401 4672 9413 4675
rect 8628 4644 9413 4672
rect 8628 4632 8634 4644
rect 9401 4641 9413 4644
rect 9447 4641 9459 4675
rect 9401 4635 9459 4641
rect 9585 4675 9643 4681
rect 9585 4641 9597 4675
rect 9631 4672 9643 4675
rect 9950 4672 9956 4684
rect 9631 4644 9956 4672
rect 9631 4641 9643 4644
rect 9585 4635 9643 4641
rect 9950 4632 9956 4644
rect 10008 4632 10014 4684
rect 10318 4632 10324 4684
rect 10376 4632 10382 4684
rect 10428 4672 10456 4712
rect 10962 4672 10968 4684
rect 10428 4644 10968 4672
rect 10962 4632 10968 4644
rect 11020 4632 11026 4684
rect 7469 4607 7527 4613
rect 4856 4576 5488 4604
rect 4856 4564 4862 4576
rect 4985 4539 5043 4545
rect 4985 4505 4997 4539
rect 5031 4505 5043 4539
rect 5460 4536 5488 4576
rect 7469 4573 7481 4607
rect 7515 4573 7527 4607
rect 7469 4567 7527 4573
rect 8389 4607 8447 4613
rect 8389 4573 8401 4607
rect 8435 4573 8447 4607
rect 8389 4567 8447 4573
rect 8941 4607 8999 4613
rect 8941 4573 8953 4607
rect 8987 4604 8999 4607
rect 9214 4604 9220 4616
rect 8987 4576 9220 4604
rect 8987 4573 8999 4576
rect 8941 4567 8999 4573
rect 9214 4564 9220 4576
rect 9272 4564 9278 4616
rect 9306 4564 9312 4616
rect 9364 4604 9370 4616
rect 9493 4607 9551 4613
rect 9493 4604 9505 4607
rect 9364 4576 9505 4604
rect 9364 4564 9370 4576
rect 9493 4573 9505 4576
rect 9539 4573 9551 4607
rect 9493 4567 9551 4573
rect 9674 4564 9680 4616
rect 9732 4564 9738 4616
rect 10042 4564 10048 4616
rect 10100 4564 10106 4616
rect 12406 4604 12434 4780
rect 12621 4607 12679 4613
rect 12621 4604 12633 4607
rect 12406 4576 12633 4604
rect 12621 4573 12633 4576
rect 12667 4604 12679 4607
rect 12986 4604 12992 4616
rect 12667 4576 12992 4604
rect 12667 4573 12679 4576
rect 12621 4567 12679 4573
rect 12986 4564 12992 4576
rect 13044 4564 13050 4616
rect 13081 4607 13139 4613
rect 13081 4573 13093 4607
rect 13127 4604 13139 4607
rect 13170 4604 13176 4616
rect 13127 4576 13176 4604
rect 13127 4573 13139 4576
rect 13081 4567 13139 4573
rect 13170 4564 13176 4576
rect 13228 4564 13234 4616
rect 5626 4536 5632 4548
rect 5460 4508 5632 4536
rect 4985 4499 5043 4505
rect 4154 4428 4160 4480
rect 4212 4428 4218 4480
rect 4614 4428 4620 4480
rect 4672 4428 4678 4480
rect 4785 4471 4843 4477
rect 4785 4437 4797 4471
rect 4831 4468 4843 4471
rect 4890 4468 4896 4480
rect 4831 4440 4896 4468
rect 4831 4437 4843 4440
rect 4785 4431 4843 4437
rect 4890 4428 4896 4440
rect 4948 4428 4954 4480
rect 5000 4468 5028 4499
rect 5626 4496 5632 4508
rect 5684 4496 5690 4548
rect 5718 4496 5724 4548
rect 5776 4496 5782 4548
rect 7377 4539 7435 4545
rect 7377 4536 7389 4539
rect 6946 4508 7389 4536
rect 7377 4505 7389 4508
rect 7423 4505 7435 4539
rect 7377 4499 7435 4505
rect 8294 4496 8300 4548
rect 8352 4536 8358 4548
rect 8573 4539 8631 4545
rect 8573 4536 8585 4539
rect 8352 4508 8585 4536
rect 8352 4496 8358 4508
rect 8573 4505 8585 4508
rect 8619 4536 8631 4539
rect 9324 4536 9352 4564
rect 10134 4536 10140 4548
rect 8619 4508 10140 4536
rect 8619 4505 8631 4508
rect 8573 4499 8631 4505
rect 10134 4496 10140 4508
rect 10192 4496 10198 4548
rect 10597 4539 10655 4545
rect 10597 4536 10609 4539
rect 10428 4508 10609 4536
rect 6086 4468 6092 4480
rect 5000 4440 6092 4468
rect 6086 4428 6092 4440
rect 6144 4428 6150 4480
rect 8662 4428 8668 4480
rect 8720 4468 8726 4480
rect 8757 4471 8815 4477
rect 8757 4468 8769 4471
rect 8720 4440 8769 4468
rect 8720 4428 8726 4440
rect 8757 4437 8769 4440
rect 8803 4437 8815 4471
rect 8757 4431 8815 4437
rect 9122 4428 9128 4480
rect 9180 4428 9186 4480
rect 9217 4471 9275 4477
rect 9217 4437 9229 4471
rect 9263 4468 9275 4471
rect 9306 4468 9312 4480
rect 9263 4440 9312 4468
rect 9263 4437 9275 4440
rect 9217 4431 9275 4437
rect 9306 4428 9312 4440
rect 9364 4428 9370 4480
rect 10229 4471 10287 4477
rect 10229 4437 10241 4471
rect 10275 4468 10287 4471
rect 10428 4468 10456 4508
rect 10597 4505 10609 4508
rect 10643 4505 10655 4539
rect 11822 4508 13124 4536
rect 10597 4499 10655 4505
rect 13096 4480 13124 4508
rect 10275 4440 10456 4468
rect 10275 4437 10287 4440
rect 10229 4431 10287 4437
rect 10778 4428 10784 4480
rect 10836 4468 10842 4480
rect 12069 4471 12127 4477
rect 12069 4468 12081 4471
rect 10836 4440 12081 4468
rect 10836 4428 10842 4440
rect 12069 4437 12081 4440
rect 12115 4437 12127 4471
rect 12069 4431 12127 4437
rect 12434 4428 12440 4480
rect 12492 4468 12498 4480
rect 12529 4471 12587 4477
rect 12529 4468 12541 4471
rect 12492 4440 12541 4468
rect 12492 4428 12498 4440
rect 12529 4437 12541 4440
rect 12575 4437 12587 4471
rect 12529 4431 12587 4437
rect 13078 4428 13084 4480
rect 13136 4428 13142 4480
rect 13262 4428 13268 4480
rect 13320 4428 13326 4480
rect 1104 4378 13708 4400
rect 1104 4326 3185 4378
rect 3237 4326 3249 4378
rect 3301 4326 3313 4378
rect 3365 4326 3377 4378
rect 3429 4326 3441 4378
rect 3493 4326 6336 4378
rect 6388 4326 6400 4378
rect 6452 4326 6464 4378
rect 6516 4326 6528 4378
rect 6580 4326 6592 4378
rect 6644 4326 9487 4378
rect 9539 4326 9551 4378
rect 9603 4326 9615 4378
rect 9667 4326 9679 4378
rect 9731 4326 9743 4378
rect 9795 4326 12638 4378
rect 12690 4326 12702 4378
rect 12754 4326 12766 4378
rect 12818 4326 12830 4378
rect 12882 4326 12894 4378
rect 12946 4326 13708 4378
rect 1104 4304 13708 4326
rect 4249 4267 4307 4273
rect 4249 4233 4261 4267
rect 4295 4264 4307 4267
rect 4338 4264 4344 4276
rect 4295 4236 4344 4264
rect 4295 4233 4307 4236
rect 4249 4227 4307 4233
rect 4338 4224 4344 4236
rect 4396 4224 4402 4276
rect 5166 4224 5172 4276
rect 5224 4264 5230 4276
rect 5534 4264 5540 4276
rect 5224 4236 5540 4264
rect 5224 4224 5230 4236
rect 5534 4224 5540 4236
rect 5592 4264 5598 4276
rect 5592 4236 5672 4264
rect 5592 4224 5598 4236
rect 5644 4205 5672 4236
rect 5718 4224 5724 4276
rect 5776 4264 5782 4276
rect 5813 4267 5871 4273
rect 5813 4264 5825 4267
rect 5776 4236 5825 4264
rect 5776 4224 5782 4236
rect 5813 4233 5825 4236
rect 5859 4233 5871 4267
rect 5813 4227 5871 4233
rect 9950 4224 9956 4276
rect 10008 4264 10014 4276
rect 10686 4264 10692 4276
rect 10008 4236 10692 4264
rect 10008 4224 10014 4236
rect 10686 4224 10692 4236
rect 10744 4264 10750 4276
rect 10781 4267 10839 4273
rect 10781 4264 10793 4267
rect 10744 4236 10793 4264
rect 10744 4224 10750 4236
rect 10781 4233 10793 4236
rect 10827 4233 10839 4267
rect 10781 4227 10839 4233
rect 10962 4224 10968 4276
rect 11020 4224 11026 4276
rect 4065 4199 4123 4205
rect 4065 4165 4077 4199
rect 4111 4196 4123 4199
rect 5445 4199 5503 4205
rect 5445 4196 5457 4199
rect 4111 4168 4384 4196
rect 4111 4165 4123 4168
rect 4065 4159 4123 4165
rect 4356 4069 4384 4168
rect 4632 4168 5457 4196
rect 4632 4137 4660 4168
rect 5445 4165 5457 4168
rect 5491 4165 5503 4199
rect 5445 4159 5503 4165
rect 5629 4199 5687 4205
rect 5629 4165 5641 4199
rect 5675 4196 5687 4199
rect 5675 4168 6132 4196
rect 5675 4165 5687 4168
rect 5629 4159 5687 4165
rect 4617 4131 4675 4137
rect 4617 4097 4629 4131
rect 4663 4097 4675 4131
rect 4617 4091 4675 4097
rect 4801 4131 4859 4137
rect 4801 4097 4813 4131
rect 4847 4128 4859 4131
rect 5258 4128 5264 4140
rect 4847 4100 5264 4128
rect 4847 4097 4859 4100
rect 4801 4091 4859 4097
rect 5258 4088 5264 4100
rect 5316 4088 5322 4140
rect 5353 4131 5411 4137
rect 5353 4097 5365 4131
rect 5399 4097 5411 4131
rect 5353 4091 5411 4097
rect 4341 4063 4399 4069
rect 4341 4029 4353 4063
rect 4387 4029 4399 4063
rect 4341 4023 4399 4029
rect 4525 4063 4583 4069
rect 4525 4029 4537 4063
rect 4571 4029 4583 4063
rect 4525 4023 4583 4029
rect 4709 4063 4767 4069
rect 4709 4029 4721 4063
rect 4755 4060 4767 4063
rect 5166 4060 5172 4072
rect 4755 4032 5172 4060
rect 4755 4029 4767 4032
rect 4709 4023 4767 4029
rect 3697 3995 3755 4001
rect 3697 3961 3709 3995
rect 3743 3992 3755 3995
rect 4246 3992 4252 4004
rect 3743 3964 4252 3992
rect 3743 3961 3755 3964
rect 3697 3955 3755 3961
rect 4246 3952 4252 3964
rect 4304 3992 4310 4004
rect 4540 3992 4568 4023
rect 5166 4020 5172 4032
rect 5224 4020 5230 4072
rect 5368 4060 5396 4091
rect 5460 4072 5488 4159
rect 5994 4088 6000 4140
rect 6052 4088 6058 4140
rect 6104 4128 6132 4168
rect 6178 4156 6184 4208
rect 6236 4196 6242 4208
rect 6517 4199 6575 4205
rect 6517 4196 6529 4199
rect 6236 4168 6529 4196
rect 6236 4156 6242 4168
rect 6517 4165 6529 4168
rect 6563 4165 6575 4199
rect 6517 4159 6575 4165
rect 6733 4199 6791 4205
rect 6733 4165 6745 4199
rect 6779 4196 6791 4199
rect 6917 4199 6975 4205
rect 6917 4196 6929 4199
rect 6779 4168 6929 4196
rect 6779 4165 6791 4168
rect 6733 4159 6791 4165
rect 6917 4165 6929 4168
rect 6963 4165 6975 4199
rect 10318 4196 10324 4208
rect 6917 4159 6975 4165
rect 9784 4168 10324 4196
rect 9784 4140 9812 4168
rect 10318 4156 10324 4168
rect 10376 4156 10382 4208
rect 10410 4156 10416 4208
rect 10468 4196 10474 4208
rect 10873 4199 10931 4205
rect 10873 4196 10885 4199
rect 10468 4168 10885 4196
rect 10468 4156 10474 4168
rect 10873 4165 10885 4168
rect 10919 4165 10931 4199
rect 10873 4159 10931 4165
rect 6822 4128 6828 4140
rect 6104 4100 6828 4128
rect 6822 4088 6828 4100
rect 6880 4088 6886 4140
rect 7009 4131 7067 4137
rect 7009 4097 7021 4131
rect 7055 4097 7067 4131
rect 7009 4091 7067 4097
rect 5276 4032 5396 4060
rect 4982 3992 4988 4004
rect 4304 3964 4384 3992
rect 4540 3964 4988 3992
rect 4304 3952 4310 3964
rect 3970 3884 3976 3936
rect 4028 3924 4034 3936
rect 4065 3927 4123 3933
rect 4065 3924 4077 3927
rect 4028 3896 4077 3924
rect 4028 3884 4034 3896
rect 4065 3893 4077 3896
rect 4111 3893 4123 3927
rect 4356 3924 4384 3964
rect 4982 3952 4988 3964
rect 5040 3992 5046 4004
rect 5276 3992 5304 4032
rect 5442 4020 5448 4072
rect 5500 4060 5506 4072
rect 7024 4060 7052 4091
rect 8386 4088 8392 4140
rect 8444 4088 8450 4140
rect 9766 4088 9772 4140
rect 9824 4088 9830 4140
rect 10045 4131 10103 4137
rect 10045 4097 10057 4131
rect 10091 4128 10103 4131
rect 10505 4131 10563 4137
rect 10091 4100 10456 4128
rect 10091 4097 10103 4100
rect 10045 4091 10103 4097
rect 7650 4060 7656 4072
rect 5500 4032 7656 4060
rect 5500 4020 5506 4032
rect 7650 4020 7656 4032
rect 7708 4020 7714 4072
rect 9122 4020 9128 4072
rect 9180 4060 9186 4072
rect 9493 4063 9551 4069
rect 9493 4060 9505 4063
rect 9180 4032 9505 4060
rect 9180 4020 9186 4032
rect 9493 4029 9505 4032
rect 9539 4029 9551 4063
rect 9493 4023 9551 4029
rect 10134 4020 10140 4072
rect 10192 4020 10198 4072
rect 10428 4060 10456 4100
rect 10505 4097 10517 4131
rect 10551 4128 10563 4131
rect 10597 4131 10655 4137
rect 10597 4128 10609 4131
rect 10551 4100 10609 4128
rect 10551 4097 10563 4100
rect 10505 4091 10563 4097
rect 10597 4097 10609 4100
rect 10643 4128 10655 4131
rect 10778 4128 10784 4140
rect 10643 4100 10784 4128
rect 10643 4097 10655 4100
rect 10597 4091 10655 4097
rect 10778 4088 10784 4100
rect 10836 4088 10842 4140
rect 11146 4088 11152 4140
rect 11204 4128 11210 4140
rect 11885 4131 11943 4137
rect 11204 4100 11836 4128
rect 11204 4088 11210 4100
rect 11808 4069 11836 4100
rect 11885 4097 11897 4131
rect 11931 4128 11943 4131
rect 12253 4131 12311 4137
rect 12253 4128 12265 4131
rect 11931 4100 12265 4128
rect 11931 4097 11943 4100
rect 11885 4091 11943 4097
rect 12253 4097 12265 4100
rect 12299 4097 12311 4131
rect 12253 4091 12311 4097
rect 12986 4088 12992 4140
rect 13044 4088 13050 4140
rect 13078 4088 13084 4140
rect 13136 4088 13142 4140
rect 11793 4063 11851 4069
rect 10428 4032 11744 4060
rect 5040 3964 5304 3992
rect 5040 3952 5046 3964
rect 5626 3952 5632 4004
rect 5684 3992 5690 4004
rect 6730 3992 6736 4004
rect 5684 3964 6736 3992
rect 5684 3952 5690 3964
rect 5077 3927 5135 3933
rect 5077 3924 5089 3927
rect 4356 3896 5089 3924
rect 4065 3887 4123 3893
rect 5077 3893 5089 3896
rect 5123 3893 5135 3927
rect 5077 3887 5135 3893
rect 5994 3884 6000 3936
rect 6052 3924 6058 3936
rect 6564 3933 6592 3964
rect 6730 3952 6736 3964
rect 6788 3952 6794 4004
rect 11716 3992 11744 4032
rect 11793 4029 11805 4063
rect 11839 4029 11851 4063
rect 11793 4023 11851 4029
rect 12805 4063 12863 4069
rect 12805 4029 12817 4063
rect 12851 4060 12863 4063
rect 13170 4060 13176 4072
rect 12851 4032 13176 4060
rect 12851 4029 12863 4032
rect 12805 4023 12863 4029
rect 12526 3992 12532 4004
rect 11716 3964 12532 3992
rect 12526 3952 12532 3964
rect 12584 3992 12590 4004
rect 12820 3992 12848 4023
rect 13170 4020 13176 4032
rect 13228 4020 13234 4072
rect 12584 3964 12848 3992
rect 12584 3952 12590 3964
rect 6365 3927 6423 3933
rect 6365 3924 6377 3927
rect 6052 3896 6377 3924
rect 6052 3884 6058 3896
rect 6365 3893 6377 3896
rect 6411 3893 6423 3927
rect 6365 3887 6423 3893
rect 6549 3927 6607 3933
rect 6549 3893 6561 3927
rect 6595 3893 6607 3927
rect 6549 3887 6607 3893
rect 8021 3927 8079 3933
rect 8021 3893 8033 3927
rect 8067 3924 8079 3927
rect 8294 3924 8300 3936
rect 8067 3896 8300 3924
rect 8067 3893 8079 3896
rect 8021 3887 8079 3893
rect 8294 3884 8300 3896
rect 8352 3884 8358 3936
rect 9398 3884 9404 3936
rect 9456 3924 9462 3936
rect 9861 3927 9919 3933
rect 9861 3924 9873 3927
rect 9456 3896 9873 3924
rect 9456 3884 9462 3896
rect 9861 3893 9873 3896
rect 9907 3893 9919 3927
rect 9861 3887 9919 3893
rect 9950 3884 9956 3936
rect 10008 3924 10014 3936
rect 10045 3927 10103 3933
rect 10045 3924 10057 3927
rect 10008 3896 10057 3924
rect 10008 3884 10014 3896
rect 10045 3893 10057 3896
rect 10091 3893 10103 3927
rect 10045 3887 10103 3893
rect 11146 3884 11152 3936
rect 11204 3884 11210 3936
rect 11514 3884 11520 3936
rect 11572 3884 11578 3936
rect 1104 3834 13708 3856
rect 1104 3782 2525 3834
rect 2577 3782 2589 3834
rect 2641 3782 2653 3834
rect 2705 3782 2717 3834
rect 2769 3782 2781 3834
rect 2833 3782 5676 3834
rect 5728 3782 5740 3834
rect 5792 3782 5804 3834
rect 5856 3782 5868 3834
rect 5920 3782 5932 3834
rect 5984 3782 8827 3834
rect 8879 3782 8891 3834
rect 8943 3782 8955 3834
rect 9007 3782 9019 3834
rect 9071 3782 9083 3834
rect 9135 3782 11978 3834
rect 12030 3782 12042 3834
rect 12094 3782 12106 3834
rect 12158 3782 12170 3834
rect 12222 3782 12234 3834
rect 12286 3782 13708 3834
rect 1104 3760 13708 3782
rect 4614 3720 4620 3732
rect 3160 3692 4620 3720
rect 842 3612 848 3664
rect 900 3652 906 3664
rect 1397 3655 1455 3661
rect 1397 3652 1409 3655
rect 900 3624 1409 3652
rect 900 3612 906 3624
rect 1397 3621 1409 3624
rect 1443 3621 1455 3655
rect 1397 3615 1455 3621
rect 3160 3525 3188 3692
rect 4614 3680 4620 3692
rect 4672 3680 4678 3732
rect 5258 3680 5264 3732
rect 5316 3720 5322 3732
rect 5537 3723 5595 3729
rect 5537 3720 5549 3723
rect 5316 3692 5549 3720
rect 5316 3680 5322 3692
rect 5537 3689 5549 3692
rect 5583 3689 5595 3723
rect 5537 3683 5595 3689
rect 7650 3680 7656 3732
rect 7708 3680 7714 3732
rect 8665 3723 8723 3729
rect 8665 3689 8677 3723
rect 8711 3720 8723 3723
rect 9198 3723 9256 3729
rect 9198 3720 9210 3723
rect 8711 3692 9210 3720
rect 8711 3689 8723 3692
rect 8665 3683 8723 3689
rect 9198 3689 9210 3692
rect 9244 3689 9256 3723
rect 9198 3683 9256 3689
rect 10686 3680 10692 3732
rect 10744 3680 10750 3732
rect 12526 3680 12532 3732
rect 12584 3680 12590 3732
rect 3510 3544 3516 3596
rect 3568 3584 3574 3596
rect 3789 3587 3847 3593
rect 3789 3584 3801 3587
rect 3568 3556 3801 3584
rect 3568 3544 3574 3556
rect 3789 3553 3801 3556
rect 3835 3584 3847 3587
rect 4062 3584 4068 3596
rect 3835 3556 4068 3584
rect 3835 3553 3847 3556
rect 3789 3547 3847 3553
rect 4062 3544 4068 3556
rect 4120 3544 4126 3596
rect 5534 3544 5540 3596
rect 5592 3584 5598 3596
rect 5905 3587 5963 3593
rect 5905 3584 5917 3587
rect 5592 3556 5917 3584
rect 5592 3544 5598 3556
rect 5905 3553 5917 3556
rect 5951 3553 5963 3587
rect 5905 3547 5963 3553
rect 8478 3544 8484 3596
rect 8536 3544 8542 3596
rect 8941 3587 8999 3593
rect 8941 3553 8953 3587
rect 8987 3584 8999 3587
rect 9766 3584 9772 3596
rect 8987 3556 9772 3584
rect 8987 3553 8999 3556
rect 8941 3547 8999 3553
rect 9766 3544 9772 3556
rect 9824 3584 9830 3596
rect 10781 3587 10839 3593
rect 10781 3584 10793 3587
rect 9824 3556 10793 3584
rect 9824 3544 9830 3556
rect 10781 3553 10793 3556
rect 10827 3553 10839 3587
rect 10781 3547 10839 3553
rect 11057 3587 11115 3593
rect 11057 3553 11069 3587
rect 11103 3584 11115 3587
rect 11514 3584 11520 3596
rect 11103 3556 11520 3584
rect 11103 3553 11115 3556
rect 11057 3547 11115 3553
rect 11514 3544 11520 3556
rect 11572 3544 11578 3596
rect 3145 3519 3203 3525
rect 3145 3485 3157 3519
rect 3191 3485 3203 3519
rect 3145 3479 3203 3485
rect 3421 3519 3479 3525
rect 3421 3485 3433 3519
rect 3467 3516 3479 3519
rect 3602 3516 3608 3528
rect 3467 3488 3608 3516
rect 3467 3485 3479 3488
rect 3421 3479 3479 3485
rect 3602 3476 3608 3488
rect 3660 3476 3666 3528
rect 5629 3519 5687 3525
rect 5629 3485 5641 3519
rect 5675 3516 5687 3519
rect 5810 3516 5816 3528
rect 5675 3488 5816 3516
rect 5675 3485 5687 3488
rect 5629 3479 5687 3485
rect 5810 3476 5816 3488
rect 5868 3476 5874 3528
rect 7926 3476 7932 3528
rect 7984 3476 7990 3528
rect 8389 3519 8447 3525
rect 8389 3485 8401 3519
rect 8435 3516 8447 3519
rect 8570 3516 8576 3528
rect 8435 3488 8576 3516
rect 8435 3485 8447 3488
rect 8389 3479 8447 3485
rect 8570 3476 8576 3488
rect 8628 3476 8634 3528
rect 13354 3476 13360 3528
rect 13412 3476 13418 3528
rect 4062 3408 4068 3460
rect 4120 3408 4126 3460
rect 6181 3451 6239 3457
rect 6181 3448 6193 3451
rect 4172 3420 4554 3448
rect 5828 3420 6193 3448
rect 3050 3340 3056 3392
rect 3108 3380 3114 3392
rect 3329 3383 3387 3389
rect 3329 3380 3341 3383
rect 3108 3352 3341 3380
rect 3108 3340 3114 3352
rect 3329 3349 3341 3352
rect 3375 3349 3387 3383
rect 3329 3343 3387 3349
rect 3513 3383 3571 3389
rect 3513 3349 3525 3383
rect 3559 3380 3571 3383
rect 4172 3380 4200 3420
rect 5828 3389 5856 3420
rect 6181 3417 6193 3420
rect 6227 3417 6239 3451
rect 6181 3411 6239 3417
rect 6914 3408 6920 3460
rect 6972 3408 6978 3460
rect 8021 3451 8079 3457
rect 8021 3417 8033 3451
rect 8067 3448 8079 3451
rect 12434 3448 12440 3460
rect 8067 3420 9706 3448
rect 12282 3420 12440 3448
rect 8067 3417 8079 3420
rect 8021 3411 8079 3417
rect 12434 3408 12440 3420
rect 12492 3408 12498 3460
rect 3559 3352 4200 3380
rect 5813 3383 5871 3389
rect 3559 3349 3571 3352
rect 3513 3343 3571 3349
rect 5813 3349 5825 3383
rect 5859 3349 5871 3383
rect 5813 3343 5871 3349
rect 1104 3290 13708 3312
rect 1104 3238 3185 3290
rect 3237 3238 3249 3290
rect 3301 3238 3313 3290
rect 3365 3238 3377 3290
rect 3429 3238 3441 3290
rect 3493 3238 6336 3290
rect 6388 3238 6400 3290
rect 6452 3238 6464 3290
rect 6516 3238 6528 3290
rect 6580 3238 6592 3290
rect 6644 3238 9487 3290
rect 9539 3238 9551 3290
rect 9603 3238 9615 3290
rect 9667 3238 9679 3290
rect 9731 3238 9743 3290
rect 9795 3238 12638 3290
rect 12690 3238 12702 3290
rect 12754 3238 12766 3290
rect 12818 3238 12830 3290
rect 12882 3238 12894 3290
rect 12946 3238 13708 3290
rect 1104 3216 13708 3238
rect 4890 3136 4896 3188
rect 4948 3176 4954 3188
rect 4985 3179 5043 3185
rect 4985 3176 4997 3179
rect 4948 3148 4997 3176
rect 4948 3136 4954 3148
rect 4985 3145 4997 3148
rect 5031 3145 5043 3179
rect 4985 3139 5043 3145
rect 5166 3136 5172 3188
rect 5224 3176 5230 3188
rect 5353 3179 5411 3185
rect 5353 3176 5365 3179
rect 5224 3148 5365 3176
rect 5224 3136 5230 3148
rect 5353 3145 5365 3148
rect 5399 3145 5411 3179
rect 5353 3139 5411 3145
rect 5813 3179 5871 3185
rect 5813 3145 5825 3179
rect 5859 3176 5871 3179
rect 6086 3176 6092 3188
rect 5859 3148 6092 3176
rect 5859 3145 5871 3148
rect 5813 3139 5871 3145
rect 6086 3136 6092 3148
rect 6144 3136 6150 3188
rect 6178 3136 6184 3188
rect 6236 3176 6242 3188
rect 6365 3179 6423 3185
rect 6365 3176 6377 3179
rect 6236 3148 6377 3176
rect 6236 3136 6242 3148
rect 6365 3145 6377 3148
rect 6411 3145 6423 3179
rect 6365 3139 6423 3145
rect 6914 3136 6920 3188
rect 6972 3176 6978 3188
rect 7009 3179 7067 3185
rect 7009 3176 7021 3179
rect 6972 3148 7021 3176
rect 6972 3136 6978 3148
rect 7009 3145 7021 3148
rect 7055 3145 7067 3179
rect 7009 3139 7067 3145
rect 8297 3179 8355 3185
rect 8297 3145 8309 3179
rect 8343 3176 8355 3179
rect 8386 3176 8392 3188
rect 8343 3148 8392 3176
rect 8343 3145 8355 3148
rect 8297 3139 8355 3145
rect 8386 3136 8392 3148
rect 8444 3136 8450 3188
rect 8662 3136 8668 3188
rect 8720 3185 8726 3188
rect 8720 3179 8739 3185
rect 8727 3145 8739 3179
rect 8720 3139 8739 3145
rect 8849 3179 8907 3185
rect 8849 3145 8861 3179
rect 8895 3176 8907 3179
rect 9214 3176 9220 3188
rect 8895 3148 9220 3176
rect 8895 3145 8907 3148
rect 8849 3139 8907 3145
rect 8720 3136 8726 3139
rect 9214 3136 9220 3148
rect 9272 3136 9278 3188
rect 9309 3179 9367 3185
rect 9309 3145 9321 3179
rect 9355 3176 9367 3179
rect 9398 3176 9404 3188
rect 9355 3148 9404 3176
rect 9355 3145 9367 3148
rect 9309 3139 9367 3145
rect 9398 3136 9404 3148
rect 9456 3136 9462 3188
rect 9493 3179 9551 3185
rect 9493 3145 9505 3179
rect 9539 3176 9551 3179
rect 10042 3176 10048 3188
rect 9539 3148 10048 3176
rect 9539 3145 9551 3148
rect 9493 3139 9551 3145
rect 10042 3136 10048 3148
rect 10100 3136 10106 3188
rect 3510 3108 3516 3120
rect 3160 3080 3516 3108
rect 3160 3049 3188 3080
rect 3510 3068 3516 3080
rect 3568 3068 3574 3120
rect 4154 3068 4160 3120
rect 4212 3068 4218 3120
rect 5537 3111 5595 3117
rect 5537 3108 5549 3111
rect 5184 3080 5549 3108
rect 5184 3049 5212 3080
rect 5537 3077 5549 3080
rect 5583 3077 5595 3111
rect 6733 3111 6791 3117
rect 6733 3108 6745 3111
rect 5537 3071 5595 3077
rect 5736 3080 6745 3108
rect 3145 3043 3203 3049
rect 3145 3009 3157 3043
rect 3191 3009 3203 3043
rect 3145 3003 3203 3009
rect 5169 3043 5227 3049
rect 5169 3009 5181 3043
rect 5215 3009 5227 3043
rect 5169 3003 5227 3009
rect 842 2932 848 2984
rect 900 2972 906 2984
rect 1397 2975 1455 2981
rect 1397 2972 1409 2975
rect 900 2944 1409 2972
rect 900 2932 906 2944
rect 1397 2941 1409 2944
rect 1443 2941 1455 2975
rect 1397 2935 1455 2941
rect 3050 2932 3056 2984
rect 3108 2972 3114 2984
rect 3421 2975 3479 2981
rect 3421 2972 3433 2975
rect 3108 2944 3433 2972
rect 3108 2932 3114 2944
rect 3421 2941 3433 2944
rect 3467 2941 3479 2975
rect 3421 2935 3479 2941
rect 4893 2975 4951 2981
rect 4893 2941 4905 2975
rect 4939 2972 4951 2975
rect 4982 2972 4988 2984
rect 4939 2944 4988 2972
rect 4939 2941 4951 2944
rect 4893 2935 4951 2941
rect 4982 2932 4988 2944
rect 5040 2972 5046 2984
rect 5184 2972 5212 3003
rect 5442 3000 5448 3052
rect 5500 3040 5506 3052
rect 5736 3049 5764 3080
rect 6733 3077 6745 3080
rect 6779 3077 6791 3111
rect 6733 3071 6791 3077
rect 8478 3068 8484 3120
rect 8536 3068 8542 3120
rect 5721 3043 5779 3049
rect 5721 3040 5733 3043
rect 5500 3012 5733 3040
rect 5500 3000 5506 3012
rect 5721 3009 5733 3012
rect 5767 3009 5779 3043
rect 5721 3003 5779 3009
rect 5813 3043 5871 3049
rect 5813 3009 5825 3043
rect 5859 3040 5871 3043
rect 6549 3043 6607 3049
rect 6549 3040 6561 3043
rect 5859 3012 6561 3040
rect 5859 3009 5871 3012
rect 5813 3003 5871 3009
rect 6549 3009 6561 3012
rect 6595 3040 6607 3043
rect 6822 3040 6828 3052
rect 6595 3012 6828 3040
rect 6595 3009 6607 3012
rect 6549 3003 6607 3009
rect 6822 3000 6828 3012
rect 6880 3000 6886 3052
rect 6917 3043 6975 3049
rect 6917 3009 6929 3043
rect 6963 3040 6975 3043
rect 7926 3040 7932 3052
rect 6963 3012 7932 3040
rect 6963 3009 6975 3012
rect 6917 3003 6975 3009
rect 7926 3000 7932 3012
rect 7984 3040 7990 3052
rect 8205 3043 8263 3049
rect 8205 3040 8217 3043
rect 7984 3012 8217 3040
rect 7984 3000 7990 3012
rect 8205 3009 8217 3012
rect 8251 3009 8263 3043
rect 8205 3003 8263 3009
rect 8570 3000 8576 3052
rect 8628 3040 8634 3052
rect 9585 3043 9643 3049
rect 9585 3040 9597 3043
rect 8628 3012 9597 3040
rect 8628 3000 8634 3012
rect 9585 3009 9597 3012
rect 9631 3009 9643 3043
rect 11146 3040 11152 3052
rect 9585 3003 9643 3009
rect 10060 3012 11152 3040
rect 5040 2944 5212 2972
rect 8941 2975 8999 2981
rect 5040 2932 5046 2944
rect 8941 2941 8953 2975
rect 8987 2972 8999 2975
rect 10060 2972 10088 3012
rect 11146 3000 11152 3012
rect 11204 3000 11210 3052
rect 8987 2944 10088 2972
rect 8987 2941 8999 2944
rect 8941 2935 8999 2941
rect 10226 2932 10232 2984
rect 10284 2972 10290 2984
rect 10686 2972 10692 2984
rect 10284 2944 10692 2972
rect 10284 2932 10290 2944
rect 10686 2932 10692 2944
rect 10744 2932 10750 2984
rect 13354 2932 13360 2984
rect 13412 2932 13418 2984
rect 9398 2904 9404 2916
rect 9232 2876 9404 2904
rect 8665 2839 8723 2845
rect 8665 2805 8677 2839
rect 8711 2836 8723 2839
rect 9232 2836 9260 2876
rect 9398 2864 9404 2876
rect 9456 2864 9462 2916
rect 8711 2808 9260 2836
rect 8711 2805 8723 2808
rect 8665 2799 8723 2805
rect 9306 2796 9312 2848
rect 9364 2796 9370 2848
rect 1104 2746 13708 2768
rect 1104 2694 2525 2746
rect 2577 2694 2589 2746
rect 2641 2694 2653 2746
rect 2705 2694 2717 2746
rect 2769 2694 2781 2746
rect 2833 2694 5676 2746
rect 5728 2694 5740 2746
rect 5792 2694 5804 2746
rect 5856 2694 5868 2746
rect 5920 2694 5932 2746
rect 5984 2694 8827 2746
rect 8879 2694 8891 2746
rect 8943 2694 8955 2746
rect 9007 2694 9019 2746
rect 9071 2694 9083 2746
rect 9135 2694 11978 2746
rect 12030 2694 12042 2746
rect 12094 2694 12106 2746
rect 12158 2694 12170 2746
rect 12222 2694 12234 2746
rect 12286 2694 13708 2746
rect 1104 2672 13708 2694
rect 4154 2592 4160 2644
rect 4212 2592 4218 2644
rect 7374 2592 7380 2644
rect 7432 2592 7438 2644
rect 10134 2496 10140 2508
rect 9416 2468 10140 2496
rect 3602 2388 3608 2440
rect 3660 2428 3666 2440
rect 4065 2431 4123 2437
rect 4065 2428 4077 2431
rect 3660 2400 4077 2428
rect 3660 2388 3666 2400
rect 4065 2397 4077 2400
rect 4111 2397 4123 2431
rect 4065 2391 4123 2397
rect 7098 2388 7104 2440
rect 7156 2428 7162 2440
rect 9416 2437 9444 2468
rect 10134 2456 10140 2468
rect 10192 2456 10198 2508
rect 7193 2431 7251 2437
rect 7193 2428 7205 2431
rect 7156 2400 7205 2428
rect 7156 2388 7162 2400
rect 7193 2397 7205 2400
rect 7239 2397 7251 2431
rect 7193 2391 7251 2397
rect 9401 2431 9459 2437
rect 9401 2397 9413 2431
rect 9447 2397 9459 2431
rect 9401 2391 9459 2397
rect 10045 2431 10103 2437
rect 10045 2397 10057 2431
rect 10091 2428 10103 2431
rect 10226 2428 10232 2440
rect 10091 2400 10232 2428
rect 10091 2397 10103 2400
rect 10045 2391 10103 2397
rect 10226 2388 10232 2400
rect 10284 2388 10290 2440
rect 10689 2431 10747 2437
rect 10689 2397 10701 2431
rect 10735 2428 10747 2431
rect 10778 2428 10784 2440
rect 10735 2400 10784 2428
rect 10735 2397 10747 2400
rect 10689 2391 10747 2397
rect 10778 2388 10784 2400
rect 10836 2388 10842 2440
rect 9030 2252 9036 2304
rect 9088 2292 9094 2304
rect 9217 2295 9275 2301
rect 9217 2292 9229 2295
rect 9088 2264 9229 2292
rect 9088 2252 9094 2264
rect 9217 2261 9229 2264
rect 9263 2261 9275 2295
rect 9217 2255 9275 2261
rect 9858 2252 9864 2304
rect 9916 2252 9922 2304
rect 10318 2252 10324 2304
rect 10376 2292 10382 2304
rect 10505 2295 10563 2301
rect 10505 2292 10517 2295
rect 10376 2264 10517 2292
rect 10376 2252 10382 2264
rect 10505 2261 10517 2264
rect 10551 2261 10563 2295
rect 10505 2255 10563 2261
rect 1104 2202 13708 2224
rect 1104 2150 3185 2202
rect 3237 2150 3249 2202
rect 3301 2150 3313 2202
rect 3365 2150 3377 2202
rect 3429 2150 3441 2202
rect 3493 2150 6336 2202
rect 6388 2150 6400 2202
rect 6452 2150 6464 2202
rect 6516 2150 6528 2202
rect 6580 2150 6592 2202
rect 6644 2150 9487 2202
rect 9539 2150 9551 2202
rect 9603 2150 9615 2202
rect 9667 2150 9679 2202
rect 9731 2150 9743 2202
rect 9795 2150 12638 2202
rect 12690 2150 12702 2202
rect 12754 2150 12766 2202
rect 12818 2150 12830 2202
rect 12882 2150 12894 2202
rect 12946 2150 13708 2202
rect 1104 2128 13708 2150
<< via1 >>
rect 2525 14662 2577 14714
rect 2589 14662 2641 14714
rect 2653 14662 2705 14714
rect 2717 14662 2769 14714
rect 2781 14662 2833 14714
rect 5676 14662 5728 14714
rect 5740 14662 5792 14714
rect 5804 14662 5856 14714
rect 5868 14662 5920 14714
rect 5932 14662 5984 14714
rect 8827 14662 8879 14714
rect 8891 14662 8943 14714
rect 8955 14662 9007 14714
rect 9019 14662 9071 14714
rect 9083 14662 9135 14714
rect 11978 14662 12030 14714
rect 12042 14662 12094 14714
rect 12106 14662 12158 14714
rect 12170 14662 12222 14714
rect 12234 14662 12286 14714
rect 3185 14118 3237 14170
rect 3249 14118 3301 14170
rect 3313 14118 3365 14170
rect 3377 14118 3429 14170
rect 3441 14118 3493 14170
rect 6336 14118 6388 14170
rect 6400 14118 6452 14170
rect 6464 14118 6516 14170
rect 6528 14118 6580 14170
rect 6592 14118 6644 14170
rect 9487 14118 9539 14170
rect 9551 14118 9603 14170
rect 9615 14118 9667 14170
rect 9679 14118 9731 14170
rect 9743 14118 9795 14170
rect 12638 14118 12690 14170
rect 12702 14118 12754 14170
rect 12766 14118 12818 14170
rect 12830 14118 12882 14170
rect 12894 14118 12946 14170
rect 9588 13948 9640 14000
rect 6460 13880 6512 13932
rect 6736 13880 6788 13932
rect 1400 13855 1452 13864
rect 1400 13821 1409 13855
rect 1409 13821 1443 13855
rect 1443 13821 1452 13855
rect 1400 13812 1452 13821
rect 5816 13855 5868 13864
rect 5816 13821 5825 13855
rect 5825 13821 5859 13855
rect 5859 13821 5868 13855
rect 5816 13812 5868 13821
rect 5540 13744 5592 13796
rect 4620 13676 4672 13728
rect 5448 13676 5500 13728
rect 9496 13855 9548 13864
rect 9496 13821 9505 13855
rect 9505 13821 9539 13855
rect 9539 13821 9548 13855
rect 9496 13812 9548 13821
rect 10232 13812 10284 13864
rect 13360 13855 13412 13864
rect 13360 13821 13369 13855
rect 13369 13821 13403 13855
rect 13403 13821 13412 13855
rect 13360 13812 13412 13821
rect 6184 13719 6236 13728
rect 6184 13685 6193 13719
rect 6193 13685 6227 13719
rect 6227 13685 6236 13719
rect 6184 13676 6236 13685
rect 6368 13719 6420 13728
rect 6368 13685 6377 13719
rect 6377 13685 6411 13719
rect 6411 13685 6420 13719
rect 6368 13676 6420 13685
rect 7932 13676 7984 13728
rect 2525 13574 2577 13626
rect 2589 13574 2641 13626
rect 2653 13574 2705 13626
rect 2717 13574 2769 13626
rect 2781 13574 2833 13626
rect 5676 13574 5728 13626
rect 5740 13574 5792 13626
rect 5804 13574 5856 13626
rect 5868 13574 5920 13626
rect 5932 13574 5984 13626
rect 8827 13574 8879 13626
rect 8891 13574 8943 13626
rect 8955 13574 9007 13626
rect 9019 13574 9071 13626
rect 9083 13574 9135 13626
rect 11978 13574 12030 13626
rect 12042 13574 12094 13626
rect 12106 13574 12158 13626
rect 12170 13574 12222 13626
rect 12234 13574 12286 13626
rect 4804 13472 4856 13524
rect 6000 13472 6052 13524
rect 6460 13472 6512 13524
rect 6828 13515 6880 13524
rect 6828 13481 6837 13515
rect 6837 13481 6871 13515
rect 6871 13481 6880 13515
rect 6828 13472 6880 13481
rect 7840 13515 7892 13524
rect 7840 13481 7849 13515
rect 7849 13481 7883 13515
rect 7883 13481 7892 13515
rect 7840 13472 7892 13481
rect 9496 13472 9548 13524
rect 9588 13515 9640 13524
rect 9588 13481 9597 13515
rect 9597 13481 9631 13515
rect 9631 13481 9640 13515
rect 9588 13472 9640 13481
rect 4160 13336 4212 13388
rect 6368 13336 6420 13388
rect 3700 13268 3752 13320
rect 4804 13311 4856 13320
rect 4804 13277 4813 13311
rect 4813 13277 4847 13311
rect 4847 13277 4856 13311
rect 4804 13268 4856 13277
rect 848 13132 900 13184
rect 2872 13132 2924 13184
rect 3516 13175 3568 13184
rect 3516 13141 3525 13175
rect 3525 13141 3559 13175
rect 3559 13141 3568 13175
rect 3516 13132 3568 13141
rect 4528 13200 4580 13252
rect 4620 13243 4672 13252
rect 4620 13209 4629 13243
rect 4629 13209 4663 13243
rect 4663 13209 4672 13243
rect 4620 13200 4672 13209
rect 7104 13311 7156 13320
rect 7104 13277 7113 13311
rect 7113 13277 7147 13311
rect 7147 13277 7156 13311
rect 7104 13268 7156 13277
rect 7196 13243 7248 13252
rect 7196 13209 7205 13243
rect 7205 13209 7239 13243
rect 7239 13209 7248 13243
rect 7196 13200 7248 13209
rect 8392 13268 8444 13320
rect 4344 13132 4396 13184
rect 5080 13132 5132 13184
rect 5540 13132 5592 13184
rect 8208 13200 8260 13252
rect 8484 13243 8536 13252
rect 8484 13209 8493 13243
rect 8493 13209 8527 13243
rect 8527 13209 8536 13243
rect 8484 13200 8536 13209
rect 9128 13311 9180 13320
rect 9128 13277 9137 13311
rect 9137 13277 9171 13311
rect 9171 13277 9180 13311
rect 9128 13268 9180 13277
rect 10416 13268 10468 13320
rect 9404 13200 9456 13252
rect 7748 13132 7800 13184
rect 8576 13175 8628 13184
rect 8576 13141 8585 13175
rect 8585 13141 8619 13175
rect 8619 13141 8628 13175
rect 8576 13132 8628 13141
rect 9864 13175 9916 13184
rect 9864 13141 9873 13175
rect 9873 13141 9907 13175
rect 9907 13141 9916 13175
rect 9864 13132 9916 13141
rect 13360 13175 13412 13184
rect 13360 13141 13369 13175
rect 13369 13141 13403 13175
rect 13403 13141 13412 13175
rect 13360 13132 13412 13141
rect 3185 13030 3237 13082
rect 3249 13030 3301 13082
rect 3313 13030 3365 13082
rect 3377 13030 3429 13082
rect 3441 13030 3493 13082
rect 6336 13030 6388 13082
rect 6400 13030 6452 13082
rect 6464 13030 6516 13082
rect 6528 13030 6580 13082
rect 6592 13030 6644 13082
rect 9487 13030 9539 13082
rect 9551 13030 9603 13082
rect 9615 13030 9667 13082
rect 9679 13030 9731 13082
rect 9743 13030 9795 13082
rect 12638 13030 12690 13082
rect 12702 13030 12754 13082
rect 12766 13030 12818 13082
rect 12830 13030 12882 13082
rect 12894 13030 12946 13082
rect 4804 12928 4856 12980
rect 5540 12928 5592 12980
rect 6092 12928 6144 12980
rect 2872 12903 2924 12912
rect 2872 12869 2881 12903
rect 2881 12869 2915 12903
rect 2915 12869 2924 12903
rect 2872 12860 2924 12869
rect 3516 12860 3568 12912
rect 7840 12971 7892 12980
rect 7840 12937 7849 12971
rect 7849 12937 7883 12971
rect 7883 12937 7892 12971
rect 7840 12928 7892 12937
rect 6000 12792 6052 12844
rect 6828 12860 6880 12912
rect 8392 12928 8444 12980
rect 8484 12928 8536 12980
rect 9128 12928 9180 12980
rect 1676 12724 1728 12776
rect 4160 12724 4212 12776
rect 4712 12767 4764 12776
rect 4712 12733 4721 12767
rect 4721 12733 4755 12767
rect 4755 12733 4764 12767
rect 4712 12724 4764 12733
rect 7104 12792 7156 12844
rect 7748 12792 7800 12844
rect 8576 12860 8628 12912
rect 9864 12860 9916 12912
rect 7932 12835 7984 12844
rect 7932 12801 7941 12835
rect 7941 12801 7975 12835
rect 7975 12801 7984 12835
rect 7932 12792 7984 12801
rect 10416 12792 10468 12844
rect 7932 12656 7984 12708
rect 6092 12588 6144 12640
rect 6828 12588 6880 12640
rect 6920 12631 6972 12640
rect 6920 12597 6929 12631
rect 6929 12597 6963 12631
rect 6963 12597 6972 12631
rect 6920 12588 6972 12597
rect 8024 12588 8076 12640
rect 8392 12588 8444 12640
rect 9404 12588 9456 12640
rect 10324 12588 10376 12640
rect 12440 12588 12492 12640
rect 2525 12486 2577 12538
rect 2589 12486 2641 12538
rect 2653 12486 2705 12538
rect 2717 12486 2769 12538
rect 2781 12486 2833 12538
rect 5676 12486 5728 12538
rect 5740 12486 5792 12538
rect 5804 12486 5856 12538
rect 5868 12486 5920 12538
rect 5932 12486 5984 12538
rect 8827 12486 8879 12538
rect 8891 12486 8943 12538
rect 8955 12486 9007 12538
rect 9019 12486 9071 12538
rect 9083 12486 9135 12538
rect 11978 12486 12030 12538
rect 12042 12486 12094 12538
rect 12106 12486 12158 12538
rect 12170 12486 12222 12538
rect 12234 12486 12286 12538
rect 4344 12427 4396 12436
rect 4344 12393 4353 12427
rect 4353 12393 4387 12427
rect 4387 12393 4396 12427
rect 4344 12384 4396 12393
rect 4712 12384 4764 12436
rect 6184 12384 6236 12436
rect 6736 12384 6788 12436
rect 8208 12427 8260 12436
rect 8208 12393 8217 12427
rect 8217 12393 8251 12427
rect 8251 12393 8260 12427
rect 8208 12384 8260 12393
rect 4620 12316 4672 12368
rect 5448 12316 5500 12368
rect 5080 12223 5132 12232
rect 5080 12189 5089 12223
rect 5089 12189 5123 12223
rect 5123 12189 5132 12223
rect 5080 12180 5132 12189
rect 5172 12223 5224 12232
rect 5172 12189 5181 12223
rect 5181 12189 5215 12223
rect 5215 12189 5224 12223
rect 5172 12180 5224 12189
rect 5448 12223 5500 12232
rect 5448 12189 5457 12223
rect 5457 12189 5491 12223
rect 5491 12189 5500 12223
rect 5448 12180 5500 12189
rect 6092 12248 6144 12300
rect 7932 12248 7984 12300
rect 10232 12248 10284 12300
rect 11520 12248 11572 12300
rect 8392 12223 8444 12232
rect 8392 12189 8401 12223
rect 8401 12189 8435 12223
rect 8435 12189 8444 12223
rect 8392 12180 8444 12189
rect 8576 12180 8628 12232
rect 5908 12155 5960 12164
rect 5908 12121 5917 12155
rect 5917 12121 5951 12155
rect 5951 12121 5960 12155
rect 5908 12112 5960 12121
rect 4160 12044 4212 12096
rect 4528 12044 4580 12096
rect 6920 12112 6972 12164
rect 9864 12112 9916 12164
rect 10324 12112 10376 12164
rect 11428 12155 11480 12164
rect 11428 12121 11437 12155
rect 11437 12121 11471 12155
rect 11471 12121 11480 12155
rect 11428 12112 11480 12121
rect 12440 12112 12492 12164
rect 6184 12044 6236 12096
rect 7196 12044 7248 12096
rect 9404 12044 9456 12096
rect 10876 12044 10928 12096
rect 12992 12044 13044 12096
rect 3185 11942 3237 11994
rect 3249 11942 3301 11994
rect 3313 11942 3365 11994
rect 3377 11942 3429 11994
rect 3441 11942 3493 11994
rect 6336 11942 6388 11994
rect 6400 11942 6452 11994
rect 6464 11942 6516 11994
rect 6528 11942 6580 11994
rect 6592 11942 6644 11994
rect 9487 11942 9539 11994
rect 9551 11942 9603 11994
rect 9615 11942 9667 11994
rect 9679 11942 9731 11994
rect 9743 11942 9795 11994
rect 12638 11942 12690 11994
rect 12702 11942 12754 11994
rect 12766 11942 12818 11994
rect 12830 11942 12882 11994
rect 12894 11942 12946 11994
rect 1676 11840 1728 11892
rect 4252 11840 4304 11892
rect 10232 11883 10284 11892
rect 10232 11849 10241 11883
rect 10241 11849 10275 11883
rect 10275 11849 10284 11883
rect 10232 11840 10284 11849
rect 10784 11840 10836 11892
rect 5172 11772 5224 11824
rect 6184 11815 6236 11824
rect 6184 11781 6193 11815
rect 6193 11781 6227 11815
rect 6227 11781 6236 11815
rect 6184 11772 6236 11781
rect 3700 11747 3752 11756
rect 3700 11713 3709 11747
rect 3709 11713 3743 11747
rect 3743 11713 3752 11747
rect 3700 11704 3752 11713
rect 8300 11772 8352 11824
rect 10968 11772 11020 11824
rect 1676 11679 1728 11688
rect 1676 11645 1685 11679
rect 1685 11645 1719 11679
rect 1719 11645 1728 11679
rect 1676 11636 1728 11645
rect 1952 11679 2004 11688
rect 1952 11645 1961 11679
rect 1961 11645 1995 11679
rect 1995 11645 2004 11679
rect 1952 11636 2004 11645
rect 5540 11636 5592 11688
rect 6552 11747 6604 11756
rect 6552 11713 6561 11747
rect 6561 11713 6595 11747
rect 6595 11713 6604 11747
rect 6552 11704 6604 11713
rect 3700 11568 3752 11620
rect 7104 11704 7156 11756
rect 11060 11747 11112 11756
rect 11060 11713 11069 11747
rect 11069 11713 11103 11747
rect 11103 11713 11112 11747
rect 11060 11704 11112 11713
rect 11428 11840 11480 11892
rect 11704 11747 11756 11756
rect 11704 11713 11713 11747
rect 11713 11713 11747 11747
rect 11747 11713 11756 11747
rect 11704 11704 11756 11713
rect 10600 11636 10652 11688
rect 12348 11704 12400 11756
rect 3792 11500 3844 11552
rect 4252 11543 4304 11552
rect 4252 11509 4261 11543
rect 4261 11509 4295 11543
rect 4295 11509 4304 11543
rect 4252 11500 4304 11509
rect 4896 11500 4948 11552
rect 6920 11543 6972 11552
rect 6920 11509 6929 11543
rect 6929 11509 6963 11543
rect 6963 11509 6972 11543
rect 6920 11500 6972 11509
rect 2525 11398 2577 11450
rect 2589 11398 2641 11450
rect 2653 11398 2705 11450
rect 2717 11398 2769 11450
rect 2781 11398 2833 11450
rect 5676 11398 5728 11450
rect 5740 11398 5792 11450
rect 5804 11398 5856 11450
rect 5868 11398 5920 11450
rect 5932 11398 5984 11450
rect 8827 11398 8879 11450
rect 8891 11398 8943 11450
rect 8955 11398 9007 11450
rect 9019 11398 9071 11450
rect 9083 11398 9135 11450
rect 11978 11398 12030 11450
rect 12042 11398 12094 11450
rect 12106 11398 12158 11450
rect 12170 11398 12222 11450
rect 12234 11398 12286 11450
rect 1952 11296 2004 11348
rect 5172 11296 5224 11348
rect 5908 11296 5960 11348
rect 6552 11296 6604 11348
rect 9404 11296 9456 11348
rect 9864 11296 9916 11348
rect 11704 11296 11756 11348
rect 12348 11339 12400 11348
rect 12348 11305 12357 11339
rect 12357 11305 12391 11339
rect 12391 11305 12400 11339
rect 12348 11296 12400 11305
rect 10968 11228 11020 11280
rect 2964 11092 3016 11144
rect 4160 11092 4212 11144
rect 4620 11135 4672 11144
rect 4620 11101 4637 11135
rect 4637 11101 4671 11135
rect 4671 11101 4672 11135
rect 4620 11092 4672 11101
rect 4896 11135 4948 11144
rect 4896 11101 4905 11135
rect 4905 11101 4939 11135
rect 4939 11101 4948 11135
rect 4896 11092 4948 11101
rect 5172 11135 5224 11144
rect 5172 11101 5181 11135
rect 5181 11101 5215 11135
rect 5215 11101 5224 11135
rect 5172 11092 5224 11101
rect 6920 11092 6972 11144
rect 8208 11092 8260 11144
rect 2412 10956 2464 11008
rect 2872 10999 2924 11008
rect 2872 10965 2881 10999
rect 2881 10965 2915 10999
rect 2915 10965 2924 10999
rect 2872 10956 2924 10965
rect 4252 11024 4304 11076
rect 7932 11024 7984 11076
rect 9220 11024 9272 11076
rect 10508 11135 10560 11144
rect 10508 11101 10517 11135
rect 10517 11101 10551 11135
rect 10551 11101 10560 11135
rect 10508 11092 10560 11101
rect 10600 11135 10652 11144
rect 10600 11101 10609 11135
rect 10609 11101 10643 11135
rect 10643 11101 10652 11135
rect 10600 11092 10652 11101
rect 10784 11135 10836 11144
rect 10784 11101 10793 11135
rect 10793 11101 10827 11135
rect 10827 11101 10836 11135
rect 10784 11092 10836 11101
rect 10876 11135 10928 11144
rect 10876 11101 10885 11135
rect 10885 11101 10919 11135
rect 10919 11101 10928 11135
rect 10876 11092 10928 11101
rect 11428 11203 11480 11212
rect 11428 11169 11437 11203
rect 11437 11169 11471 11203
rect 11471 11169 11480 11203
rect 11428 11160 11480 11169
rect 11612 11203 11664 11212
rect 11612 11169 11620 11203
rect 11620 11169 11654 11203
rect 11654 11169 11664 11203
rect 11612 11160 11664 11169
rect 11060 11024 11112 11076
rect 11796 11092 11848 11144
rect 12256 11228 12308 11280
rect 12072 11160 12124 11212
rect 12256 11135 12308 11144
rect 12256 11101 12265 11135
rect 12265 11101 12299 11135
rect 12299 11101 12308 11135
rect 12256 11092 12308 11101
rect 12992 11160 13044 11212
rect 12072 11024 12124 11076
rect 12348 11024 12400 11076
rect 4528 10956 4580 11008
rect 4620 10956 4672 11008
rect 5448 10956 5500 11008
rect 8392 10956 8444 11008
rect 9956 10956 10008 11008
rect 11152 10956 11204 11008
rect 12256 10956 12308 11008
rect 12532 10956 12584 11008
rect 3185 10854 3237 10906
rect 3249 10854 3301 10906
rect 3313 10854 3365 10906
rect 3377 10854 3429 10906
rect 3441 10854 3493 10906
rect 6336 10854 6388 10906
rect 6400 10854 6452 10906
rect 6464 10854 6516 10906
rect 6528 10854 6580 10906
rect 6592 10854 6644 10906
rect 9487 10854 9539 10906
rect 9551 10854 9603 10906
rect 9615 10854 9667 10906
rect 9679 10854 9731 10906
rect 9743 10854 9795 10906
rect 12638 10854 12690 10906
rect 12702 10854 12754 10906
rect 12766 10854 12818 10906
rect 12830 10854 12882 10906
rect 12894 10854 12946 10906
rect 4160 10752 4212 10804
rect 3056 10684 3108 10736
rect 3792 10727 3844 10736
rect 3792 10693 3801 10727
rect 3801 10693 3835 10727
rect 3835 10693 3844 10727
rect 3792 10684 3844 10693
rect 1492 10659 1544 10668
rect 1492 10625 1501 10659
rect 1501 10625 1535 10659
rect 1535 10625 1544 10659
rect 1492 10616 1544 10625
rect 4160 10616 4212 10668
rect 5540 10752 5592 10804
rect 8392 10752 8444 10804
rect 9404 10752 9456 10804
rect 9588 10752 9640 10804
rect 5908 10727 5960 10736
rect 5908 10693 5917 10727
rect 5917 10693 5951 10727
rect 5951 10693 5960 10727
rect 5908 10684 5960 10693
rect 5264 10659 5316 10668
rect 5264 10625 5273 10659
rect 5273 10625 5307 10659
rect 5307 10625 5316 10659
rect 5264 10616 5316 10625
rect 5356 10659 5408 10668
rect 5356 10625 5365 10659
rect 5365 10625 5399 10659
rect 5399 10625 5408 10659
rect 5356 10616 5408 10625
rect 6736 10616 6788 10668
rect 9680 10684 9732 10736
rect 10876 10752 10928 10804
rect 11428 10752 11480 10804
rect 11704 10752 11756 10804
rect 10600 10684 10652 10736
rect 1676 10548 1728 10600
rect 3424 10412 3476 10464
rect 4528 10548 4580 10600
rect 4804 10548 4856 10600
rect 5908 10548 5960 10600
rect 6828 10548 6880 10600
rect 8116 10616 8168 10668
rect 8576 10616 8628 10668
rect 9312 10616 9364 10668
rect 4436 10480 4488 10532
rect 4712 10480 4764 10532
rect 4344 10412 4396 10464
rect 5356 10480 5408 10532
rect 9496 10591 9548 10600
rect 9496 10557 9505 10591
rect 9505 10557 9539 10591
rect 9539 10557 9548 10591
rect 9496 10548 9548 10557
rect 9588 10591 9640 10600
rect 9588 10557 9597 10591
rect 9597 10557 9631 10591
rect 9631 10557 9640 10591
rect 9588 10548 9640 10557
rect 9956 10616 10008 10668
rect 10324 10616 10376 10668
rect 10784 10616 10836 10668
rect 12532 10684 12584 10736
rect 11152 10616 11204 10668
rect 11520 10659 11572 10668
rect 11520 10625 11529 10659
rect 11529 10625 11563 10659
rect 11563 10625 11572 10659
rect 11520 10616 11572 10625
rect 7840 10480 7892 10532
rect 8484 10480 8536 10532
rect 9220 10480 9272 10532
rect 8116 10412 8168 10464
rect 8208 10455 8260 10464
rect 8208 10421 8217 10455
rect 8217 10421 8251 10455
rect 8251 10421 8260 10455
rect 8208 10412 8260 10421
rect 8576 10412 8628 10464
rect 11244 10548 11296 10600
rect 11060 10412 11112 10464
rect 12256 10412 12308 10464
rect 12348 10412 12400 10464
rect 2525 10310 2577 10362
rect 2589 10310 2641 10362
rect 2653 10310 2705 10362
rect 2717 10310 2769 10362
rect 2781 10310 2833 10362
rect 5676 10310 5728 10362
rect 5740 10310 5792 10362
rect 5804 10310 5856 10362
rect 5868 10310 5920 10362
rect 5932 10310 5984 10362
rect 8827 10310 8879 10362
rect 8891 10310 8943 10362
rect 8955 10310 9007 10362
rect 9019 10310 9071 10362
rect 9083 10310 9135 10362
rect 11978 10310 12030 10362
rect 12042 10310 12094 10362
rect 12106 10310 12158 10362
rect 12170 10310 12222 10362
rect 12234 10310 12286 10362
rect 1492 10208 1544 10260
rect 2964 10208 3016 10260
rect 3332 10208 3384 10260
rect 3792 10208 3844 10260
rect 4712 10208 4764 10260
rect 2412 10004 2464 10056
rect 3332 10047 3384 10056
rect 3332 10013 3341 10047
rect 3341 10013 3375 10047
rect 3375 10013 3384 10047
rect 3332 10004 3384 10013
rect 3424 10047 3476 10056
rect 3424 10013 3433 10047
rect 3433 10013 3467 10047
rect 3467 10013 3476 10047
rect 3424 10004 3476 10013
rect 4252 10072 4304 10124
rect 2872 9868 2924 9920
rect 2964 9868 3016 9920
rect 4344 10047 4396 10056
rect 4344 10013 4353 10047
rect 4353 10013 4387 10047
rect 4387 10013 4396 10047
rect 4344 10004 4396 10013
rect 4436 10047 4488 10056
rect 4436 10013 4445 10047
rect 4445 10013 4479 10047
rect 4479 10013 4488 10047
rect 4436 10004 4488 10013
rect 9404 10208 9456 10260
rect 8392 10140 8444 10192
rect 5172 10072 5224 10124
rect 7104 10004 7156 10056
rect 4620 9936 4672 9988
rect 4068 9868 4120 9920
rect 4160 9868 4212 9920
rect 5356 9868 5408 9920
rect 8208 10004 8260 10056
rect 8484 10047 8536 10056
rect 8484 10013 8493 10047
rect 8493 10013 8527 10047
rect 8527 10013 8536 10047
rect 8484 10004 8536 10013
rect 9680 10140 9732 10192
rect 11244 10208 11296 10260
rect 9956 10072 10008 10124
rect 11796 10140 11848 10192
rect 11888 10072 11940 10124
rect 12532 10072 12584 10124
rect 8116 9868 8168 9920
rect 9220 9936 9272 9988
rect 8392 9868 8444 9920
rect 8668 9868 8720 9920
rect 9312 9911 9364 9920
rect 9312 9877 9321 9911
rect 9321 9877 9355 9911
rect 9355 9877 9364 9911
rect 9312 9868 9364 9877
rect 11428 10004 11480 10056
rect 11704 10047 11756 10056
rect 11704 10013 11713 10047
rect 11713 10013 11747 10047
rect 11747 10013 11756 10047
rect 11704 10004 11756 10013
rect 12072 10047 12124 10056
rect 12072 10013 12081 10047
rect 12081 10013 12115 10047
rect 12115 10013 12124 10047
rect 12072 10004 12124 10013
rect 13268 10004 13320 10056
rect 12532 9979 12584 9988
rect 12532 9945 12541 9979
rect 12541 9945 12575 9979
rect 12575 9945 12584 9979
rect 12532 9936 12584 9945
rect 10416 9868 10468 9920
rect 11060 9868 11112 9920
rect 11336 9911 11388 9920
rect 11336 9877 11345 9911
rect 11345 9877 11379 9911
rect 11379 9877 11388 9911
rect 11336 9868 11388 9877
rect 11428 9868 11480 9920
rect 11796 9911 11848 9920
rect 11796 9877 11805 9911
rect 11805 9877 11839 9911
rect 11839 9877 11848 9911
rect 11796 9868 11848 9877
rect 11888 9868 11940 9920
rect 12348 9868 12400 9920
rect 3185 9766 3237 9818
rect 3249 9766 3301 9818
rect 3313 9766 3365 9818
rect 3377 9766 3429 9818
rect 3441 9766 3493 9818
rect 6336 9766 6388 9818
rect 6400 9766 6452 9818
rect 6464 9766 6516 9818
rect 6528 9766 6580 9818
rect 6592 9766 6644 9818
rect 9487 9766 9539 9818
rect 9551 9766 9603 9818
rect 9615 9766 9667 9818
rect 9679 9766 9731 9818
rect 9743 9766 9795 9818
rect 12638 9766 12690 9818
rect 12702 9766 12754 9818
rect 12766 9766 12818 9818
rect 12830 9766 12882 9818
rect 12894 9766 12946 9818
rect 5264 9664 5316 9716
rect 8484 9664 8536 9716
rect 9128 9664 9180 9716
rect 9956 9664 10008 9716
rect 10508 9664 10560 9716
rect 11612 9664 11664 9716
rect 12072 9664 12124 9716
rect 3056 9596 3108 9648
rect 3700 9596 3752 9648
rect 4252 9596 4304 9648
rect 5356 9596 5408 9648
rect 8116 9596 8168 9648
rect 9220 9596 9272 9648
rect 12348 9596 12400 9648
rect 2872 9460 2924 9512
rect 4160 9528 4212 9580
rect 4344 9571 4396 9580
rect 4344 9537 4353 9571
rect 4353 9537 4387 9571
rect 4387 9537 4396 9571
rect 4344 9528 4396 9537
rect 4436 9571 4488 9580
rect 4436 9537 4445 9571
rect 4445 9537 4479 9571
rect 4479 9537 4488 9571
rect 4436 9528 4488 9537
rect 4528 9460 4580 9512
rect 3884 9392 3936 9444
rect 7932 9571 7984 9580
rect 7932 9537 7941 9571
rect 7941 9537 7975 9571
rect 7975 9537 7984 9571
rect 7932 9528 7984 9537
rect 11520 9571 11572 9580
rect 11520 9537 11529 9571
rect 11529 9537 11563 9571
rect 11563 9537 11572 9571
rect 11520 9528 11572 9537
rect 11060 9460 11112 9512
rect 13268 9503 13320 9512
rect 13268 9469 13277 9503
rect 13277 9469 13311 9503
rect 13311 9469 13320 9503
rect 13268 9460 13320 9469
rect 3148 9367 3200 9376
rect 3148 9333 3157 9367
rect 3157 9333 3191 9367
rect 3191 9333 3200 9367
rect 3148 9324 3200 9333
rect 4804 9367 4856 9376
rect 4804 9333 4813 9367
rect 4813 9333 4847 9367
rect 4847 9333 4856 9367
rect 4804 9324 4856 9333
rect 5356 9324 5408 9376
rect 2525 9222 2577 9274
rect 2589 9222 2641 9274
rect 2653 9222 2705 9274
rect 2717 9222 2769 9274
rect 2781 9222 2833 9274
rect 5676 9222 5728 9274
rect 5740 9222 5792 9274
rect 5804 9222 5856 9274
rect 5868 9222 5920 9274
rect 5932 9222 5984 9274
rect 8827 9222 8879 9274
rect 8891 9222 8943 9274
rect 8955 9222 9007 9274
rect 9019 9222 9071 9274
rect 9083 9222 9135 9274
rect 11978 9222 12030 9274
rect 12042 9222 12094 9274
rect 12106 9222 12158 9274
rect 12170 9222 12222 9274
rect 12234 9222 12286 9274
rect 3148 9120 3200 9172
rect 4160 9120 4212 9172
rect 8392 9163 8444 9172
rect 8392 9129 8401 9163
rect 8401 9129 8435 9163
rect 8435 9129 8444 9163
rect 8392 9120 8444 9129
rect 8576 9163 8628 9172
rect 8576 9129 8585 9163
rect 8585 9129 8619 9163
rect 8619 9129 8628 9163
rect 8576 9120 8628 9129
rect 11060 9163 11112 9172
rect 11060 9129 11069 9163
rect 11069 9129 11103 9163
rect 11103 9129 11112 9163
rect 11060 9120 11112 9129
rect 12348 9120 12400 9172
rect 4344 9052 4396 9104
rect 5448 9052 5500 9104
rect 11336 9052 11388 9104
rect 6828 8984 6880 9036
rect 6920 8984 6972 9036
rect 8208 9027 8260 9036
rect 8208 8993 8217 9027
rect 8217 8993 8251 9027
rect 8251 8993 8260 9027
rect 8208 8984 8260 8993
rect 1952 8780 2004 8832
rect 5356 8959 5408 8968
rect 5356 8925 5365 8959
rect 5365 8925 5399 8959
rect 5399 8925 5408 8959
rect 5356 8916 5408 8925
rect 5448 8916 5500 8968
rect 2964 8891 3016 8900
rect 2964 8857 2973 8891
rect 2973 8857 3007 8891
rect 3007 8857 3016 8891
rect 2964 8848 3016 8857
rect 3884 8891 3936 8900
rect 3884 8857 3893 8891
rect 3893 8857 3927 8891
rect 3927 8857 3936 8891
rect 3884 8848 3936 8857
rect 4436 8848 4488 8900
rect 5172 8848 5224 8900
rect 6552 8959 6604 8968
rect 6552 8925 6561 8959
rect 6561 8925 6595 8959
rect 6595 8925 6604 8959
rect 6552 8916 6604 8925
rect 8576 8916 8628 8968
rect 10324 8916 10376 8968
rect 11612 9027 11664 9036
rect 11612 8993 11621 9027
rect 11621 8993 11655 9027
rect 11655 8993 11664 9027
rect 11612 8984 11664 8993
rect 13268 9027 13320 9036
rect 13268 8993 13277 9027
rect 13277 8993 13311 9027
rect 13311 8993 13320 9027
rect 13268 8984 13320 8993
rect 9404 8848 9456 8900
rect 10048 8848 10100 8900
rect 10784 8959 10836 8968
rect 10784 8925 10793 8959
rect 10793 8925 10827 8959
rect 10827 8925 10836 8959
rect 10784 8916 10836 8925
rect 11704 8848 11756 8900
rect 12348 8916 12400 8968
rect 3516 8780 3568 8832
rect 8392 8780 8444 8832
rect 3185 8678 3237 8730
rect 3249 8678 3301 8730
rect 3313 8678 3365 8730
rect 3377 8678 3429 8730
rect 3441 8678 3493 8730
rect 6336 8678 6388 8730
rect 6400 8678 6452 8730
rect 6464 8678 6516 8730
rect 6528 8678 6580 8730
rect 6592 8678 6644 8730
rect 9487 8678 9539 8730
rect 9551 8678 9603 8730
rect 9615 8678 9667 8730
rect 9679 8678 9731 8730
rect 9743 8678 9795 8730
rect 12638 8678 12690 8730
rect 12702 8678 12754 8730
rect 12766 8678 12818 8730
rect 12830 8678 12882 8730
rect 12894 8678 12946 8730
rect 1952 8551 2004 8560
rect 1952 8517 1961 8551
rect 1961 8517 1995 8551
rect 1995 8517 2004 8551
rect 1952 8508 2004 8517
rect 2964 8508 3016 8560
rect 3516 8619 3568 8628
rect 3516 8585 3525 8619
rect 3525 8585 3559 8619
rect 3559 8585 3568 8619
rect 3516 8576 3568 8585
rect 3884 8576 3936 8628
rect 6736 8576 6788 8628
rect 7656 8619 7708 8628
rect 7656 8585 7665 8619
rect 7665 8585 7699 8619
rect 7699 8585 7708 8619
rect 7656 8576 7708 8585
rect 8300 8619 8352 8628
rect 8300 8585 8309 8619
rect 8309 8585 8343 8619
rect 8343 8585 8352 8619
rect 8300 8576 8352 8585
rect 8484 8576 8536 8628
rect 8668 8576 8720 8628
rect 1676 8483 1728 8492
rect 1676 8449 1685 8483
rect 1685 8449 1719 8483
rect 1719 8449 1728 8483
rect 1676 8440 1728 8449
rect 4344 8440 4396 8492
rect 5356 8440 5408 8492
rect 6828 8483 6880 8492
rect 6828 8449 6837 8483
rect 6837 8449 6871 8483
rect 6871 8449 6880 8483
rect 7932 8508 7984 8560
rect 9220 8508 9272 8560
rect 6828 8440 6880 8449
rect 6644 8415 6696 8424
rect 6644 8381 6653 8415
rect 6653 8381 6687 8415
rect 6687 8381 6696 8415
rect 6644 8372 6696 8381
rect 7840 8372 7892 8424
rect 8392 8440 8444 8492
rect 8668 8483 8720 8492
rect 8668 8449 8677 8483
rect 8677 8449 8711 8483
rect 8711 8449 8720 8483
rect 8668 8440 8720 8449
rect 10600 8508 10652 8560
rect 11336 8508 11388 8560
rect 11888 8508 11940 8560
rect 10876 8440 10928 8492
rect 8484 8415 8536 8424
rect 8484 8381 8493 8415
rect 8493 8381 8527 8415
rect 8527 8381 8536 8415
rect 8484 8372 8536 8381
rect 4712 8236 4764 8288
rect 6736 8236 6788 8288
rect 7288 8279 7340 8288
rect 7288 8245 7297 8279
rect 7297 8245 7331 8279
rect 7331 8245 7340 8279
rect 7288 8236 7340 8245
rect 8392 8347 8444 8356
rect 8392 8313 8401 8347
rect 8401 8313 8435 8347
rect 8435 8313 8444 8347
rect 8392 8304 8444 8313
rect 8668 8236 8720 8288
rect 10140 8236 10192 8288
rect 10784 8236 10836 8288
rect 2525 8134 2577 8186
rect 2589 8134 2641 8186
rect 2653 8134 2705 8186
rect 2717 8134 2769 8186
rect 2781 8134 2833 8186
rect 5676 8134 5728 8186
rect 5740 8134 5792 8186
rect 5804 8134 5856 8186
rect 5868 8134 5920 8186
rect 5932 8134 5984 8186
rect 8827 8134 8879 8186
rect 8891 8134 8943 8186
rect 8955 8134 9007 8186
rect 9019 8134 9071 8186
rect 9083 8134 9135 8186
rect 11978 8134 12030 8186
rect 12042 8134 12094 8186
rect 12106 8134 12158 8186
rect 12170 8134 12222 8186
rect 12234 8134 12286 8186
rect 2964 8032 3016 8084
rect 4712 8075 4764 8084
rect 4712 8041 4721 8075
rect 4721 8041 4755 8075
rect 4755 8041 4764 8075
rect 4712 8032 4764 8041
rect 4344 8007 4396 8016
rect 4344 7973 4353 8007
rect 4353 7973 4387 8007
rect 4387 7973 4396 8007
rect 4344 7964 4396 7973
rect 8484 7964 8536 8016
rect 2872 7871 2924 7880
rect 2872 7837 2881 7871
rect 2881 7837 2915 7871
rect 2915 7837 2924 7871
rect 2872 7828 2924 7837
rect 5172 7871 5224 7880
rect 5172 7837 5181 7871
rect 5181 7837 5215 7871
rect 5215 7837 5224 7871
rect 5172 7828 5224 7837
rect 4436 7760 4488 7812
rect 5356 7828 5408 7880
rect 7656 7828 7708 7880
rect 8300 7828 8352 7880
rect 8760 7871 8812 7880
rect 8760 7837 8769 7871
rect 8769 7837 8803 7871
rect 8803 7837 8812 7871
rect 8760 7828 8812 7837
rect 10140 7964 10192 8016
rect 9956 7871 10008 7880
rect 9956 7837 9965 7871
rect 9965 7837 9999 7871
rect 9999 7837 10008 7871
rect 9956 7828 10008 7837
rect 10048 7828 10100 7880
rect 10600 7896 10652 7948
rect 11152 7896 11204 7948
rect 10324 7828 10376 7880
rect 10876 7871 10928 7880
rect 10876 7837 10885 7871
rect 10885 7837 10919 7871
rect 10919 7837 10928 7871
rect 10876 7828 10928 7837
rect 11060 7828 11112 7880
rect 12348 7964 12400 8016
rect 11612 7896 11664 7948
rect 11704 7871 11756 7880
rect 11704 7837 11713 7871
rect 11713 7837 11747 7871
rect 11747 7837 11756 7871
rect 11704 7828 11756 7837
rect 11796 7760 11848 7812
rect 4712 7735 4764 7744
rect 4712 7701 4721 7735
rect 4721 7701 4755 7735
rect 4755 7701 4764 7735
rect 4712 7692 4764 7701
rect 5908 7692 5960 7744
rect 7288 7692 7340 7744
rect 8484 7735 8536 7744
rect 8484 7701 8493 7735
rect 8493 7701 8527 7735
rect 8527 7701 8536 7735
rect 8484 7692 8536 7701
rect 9864 7692 9916 7744
rect 10784 7692 10836 7744
rect 11060 7692 11112 7744
rect 11244 7735 11296 7744
rect 11244 7701 11253 7735
rect 11253 7701 11287 7735
rect 11287 7701 11296 7735
rect 11244 7692 11296 7701
rect 12256 7692 12308 7744
rect 3185 7590 3237 7642
rect 3249 7590 3301 7642
rect 3313 7590 3365 7642
rect 3377 7590 3429 7642
rect 3441 7590 3493 7642
rect 6336 7590 6388 7642
rect 6400 7590 6452 7642
rect 6464 7590 6516 7642
rect 6528 7590 6580 7642
rect 6592 7590 6644 7642
rect 9487 7590 9539 7642
rect 9551 7590 9603 7642
rect 9615 7590 9667 7642
rect 9679 7590 9731 7642
rect 9743 7590 9795 7642
rect 12638 7590 12690 7642
rect 12702 7590 12754 7642
rect 12766 7590 12818 7642
rect 12830 7590 12882 7642
rect 12894 7590 12946 7642
rect 5172 7488 5224 7540
rect 2320 7148 2372 7200
rect 3516 7395 3568 7404
rect 3516 7361 3525 7395
rect 3525 7361 3559 7395
rect 3559 7361 3568 7395
rect 3516 7352 3568 7361
rect 3792 7420 3844 7472
rect 7196 7488 7248 7540
rect 8576 7488 8628 7540
rect 8852 7488 8904 7540
rect 5908 7463 5960 7472
rect 5908 7429 5917 7463
rect 5917 7429 5951 7463
rect 5951 7429 5960 7463
rect 5908 7420 5960 7429
rect 3976 7395 4028 7404
rect 3976 7361 3985 7395
rect 3985 7361 4019 7395
rect 4019 7361 4028 7395
rect 3976 7352 4028 7361
rect 6644 7420 6696 7472
rect 7104 7420 7156 7472
rect 3608 7216 3660 7268
rect 3700 7148 3752 7200
rect 6736 7352 6788 7404
rect 7380 7352 7432 7404
rect 8576 7352 8628 7404
rect 9956 7488 10008 7540
rect 11060 7488 11112 7540
rect 11704 7488 11756 7540
rect 9864 7420 9916 7472
rect 11244 7420 11296 7472
rect 9404 7352 9456 7404
rect 6184 7327 6236 7336
rect 6184 7293 6193 7327
rect 6193 7293 6227 7327
rect 6227 7293 6236 7327
rect 6184 7284 6236 7293
rect 8668 7284 8720 7336
rect 9496 7327 9548 7336
rect 9496 7293 9505 7327
rect 9505 7293 9539 7327
rect 9539 7293 9548 7327
rect 9496 7284 9548 7293
rect 10784 7284 10836 7336
rect 4620 7148 4672 7200
rect 8852 7148 8904 7200
rect 10508 7148 10560 7200
rect 11428 7352 11480 7404
rect 11612 7352 11664 7404
rect 11796 7395 11848 7404
rect 11796 7361 11805 7395
rect 11805 7361 11839 7395
rect 11839 7361 11848 7395
rect 11796 7352 11848 7361
rect 12532 7420 12584 7472
rect 11152 7284 11204 7336
rect 13268 7284 13320 7336
rect 12256 7191 12308 7200
rect 12256 7157 12265 7191
rect 12265 7157 12299 7191
rect 12299 7157 12308 7191
rect 12256 7148 12308 7157
rect 12532 7191 12584 7200
rect 12532 7157 12541 7191
rect 12541 7157 12575 7191
rect 12575 7157 12584 7191
rect 12532 7148 12584 7157
rect 12900 7191 12952 7200
rect 12900 7157 12909 7191
rect 12909 7157 12943 7191
rect 12943 7157 12952 7191
rect 12900 7148 12952 7157
rect 13176 7191 13228 7200
rect 13176 7157 13185 7191
rect 13185 7157 13219 7191
rect 13219 7157 13228 7191
rect 13176 7148 13228 7157
rect 2525 7046 2577 7098
rect 2589 7046 2641 7098
rect 2653 7046 2705 7098
rect 2717 7046 2769 7098
rect 2781 7046 2833 7098
rect 5676 7046 5728 7098
rect 5740 7046 5792 7098
rect 5804 7046 5856 7098
rect 5868 7046 5920 7098
rect 5932 7046 5984 7098
rect 8827 7046 8879 7098
rect 8891 7046 8943 7098
rect 8955 7046 9007 7098
rect 9019 7046 9071 7098
rect 9083 7046 9135 7098
rect 11978 7046 12030 7098
rect 12042 7046 12094 7098
rect 12106 7046 12158 7098
rect 12170 7046 12222 7098
rect 12234 7046 12286 7098
rect 2320 6987 2372 6996
rect 2320 6953 2329 6987
rect 2329 6953 2363 6987
rect 2363 6953 2372 6987
rect 2320 6944 2372 6953
rect 2964 6944 3016 6996
rect 2136 6919 2188 6928
rect 2136 6885 2145 6919
rect 2145 6885 2179 6919
rect 2179 6885 2188 6919
rect 2136 6876 2188 6885
rect 1860 6783 1912 6792
rect 1860 6749 1869 6783
rect 1869 6749 1903 6783
rect 1903 6749 1912 6783
rect 1860 6740 1912 6749
rect 2504 6808 2556 6860
rect 3332 6876 3384 6928
rect 3884 6876 3936 6928
rect 4436 6944 4488 6996
rect 9312 6944 9364 6996
rect 9680 6944 9732 6996
rect 10324 6944 10376 6996
rect 11244 6944 11296 6996
rect 12532 6944 12584 6996
rect 2688 6808 2740 6860
rect 3608 6808 3660 6860
rect 8300 6876 8352 6928
rect 8852 6876 8904 6928
rect 9220 6876 9272 6928
rect 10692 6876 10744 6928
rect 1492 6672 1544 6724
rect 3056 6672 3108 6724
rect 3332 6783 3384 6792
rect 3332 6749 3341 6783
rect 3341 6749 3375 6783
rect 3375 6749 3384 6783
rect 3332 6740 3384 6749
rect 3516 6740 3568 6792
rect 4068 6851 4120 6860
rect 4068 6817 4077 6851
rect 4077 6817 4111 6851
rect 4111 6817 4120 6851
rect 4068 6808 4120 6817
rect 4896 6808 4948 6860
rect 6644 6851 6696 6860
rect 6644 6817 6653 6851
rect 6653 6817 6687 6851
rect 6687 6817 6696 6851
rect 6644 6808 6696 6817
rect 9496 6808 9548 6860
rect 10416 6808 10468 6860
rect 13268 6851 13320 6860
rect 13268 6817 13277 6851
rect 13277 6817 13311 6851
rect 13311 6817 13320 6851
rect 13268 6808 13320 6817
rect 3792 6783 3844 6792
rect 3792 6749 3801 6783
rect 3801 6749 3835 6783
rect 3835 6749 3844 6783
rect 3792 6740 3844 6749
rect 3976 6783 4028 6792
rect 3976 6749 3985 6783
rect 3985 6749 4019 6783
rect 4019 6749 4028 6783
rect 3976 6740 4028 6749
rect 3516 6604 3568 6656
rect 3884 6604 3936 6656
rect 4160 6604 4212 6656
rect 4344 6715 4396 6724
rect 4344 6681 4353 6715
rect 4353 6681 4387 6715
rect 4387 6681 4396 6715
rect 4344 6672 4396 6681
rect 9220 6783 9272 6792
rect 9220 6749 9229 6783
rect 9229 6749 9263 6783
rect 9263 6749 9272 6783
rect 9220 6740 9272 6749
rect 10048 6783 10100 6792
rect 10048 6749 10057 6783
rect 10057 6749 10091 6783
rect 10091 6749 10100 6783
rect 10048 6740 10100 6749
rect 10140 6783 10192 6792
rect 10140 6749 10149 6783
rect 10149 6749 10183 6783
rect 10183 6749 10192 6783
rect 10140 6740 10192 6749
rect 10232 6740 10284 6792
rect 10784 6783 10836 6792
rect 10784 6749 10793 6783
rect 10793 6749 10827 6783
rect 10827 6749 10836 6783
rect 10784 6740 10836 6749
rect 10876 6783 10928 6792
rect 10876 6749 10885 6783
rect 10885 6749 10919 6783
rect 10919 6749 10928 6783
rect 10876 6740 10928 6749
rect 7380 6672 7432 6724
rect 8300 6672 8352 6724
rect 5816 6647 5868 6656
rect 5816 6613 5825 6647
rect 5825 6613 5859 6647
rect 5859 6613 5868 6647
rect 5816 6604 5868 6613
rect 11428 6740 11480 6792
rect 12900 6740 12952 6792
rect 11336 6672 11388 6724
rect 9036 6604 9088 6656
rect 9680 6604 9732 6656
rect 9864 6647 9916 6656
rect 9864 6613 9873 6647
rect 9873 6613 9907 6647
rect 9907 6613 9916 6647
rect 9864 6604 9916 6613
rect 10048 6604 10100 6656
rect 10600 6647 10652 6656
rect 10600 6613 10609 6647
rect 10609 6613 10643 6647
rect 10643 6613 10652 6647
rect 10600 6604 10652 6613
rect 11060 6647 11112 6656
rect 11060 6613 11069 6647
rect 11069 6613 11103 6647
rect 11103 6613 11112 6647
rect 11060 6604 11112 6613
rect 3185 6502 3237 6554
rect 3249 6502 3301 6554
rect 3313 6502 3365 6554
rect 3377 6502 3429 6554
rect 3441 6502 3493 6554
rect 6336 6502 6388 6554
rect 6400 6502 6452 6554
rect 6464 6502 6516 6554
rect 6528 6502 6580 6554
rect 6592 6502 6644 6554
rect 9487 6502 9539 6554
rect 9551 6502 9603 6554
rect 9615 6502 9667 6554
rect 9679 6502 9731 6554
rect 9743 6502 9795 6554
rect 12638 6502 12690 6554
rect 12702 6502 12754 6554
rect 12766 6502 12818 6554
rect 12830 6502 12882 6554
rect 12894 6502 12946 6554
rect 4068 6400 4120 6452
rect 4344 6400 4396 6452
rect 4712 6400 4764 6452
rect 3056 6332 3108 6384
rect 1492 6307 1544 6316
rect 1492 6273 1501 6307
rect 1501 6273 1535 6307
rect 1535 6273 1544 6307
rect 1492 6264 1544 6273
rect 1768 6307 1820 6316
rect 1768 6273 1777 6307
rect 1777 6273 1811 6307
rect 1811 6273 1820 6307
rect 1768 6264 1820 6273
rect 4528 6332 4580 6384
rect 6092 6332 6144 6384
rect 8300 6400 8352 6452
rect 9036 6400 9088 6452
rect 3884 6264 3936 6316
rect 3424 6196 3476 6248
rect 4160 6307 4212 6316
rect 4160 6273 4169 6307
rect 4169 6273 4203 6307
rect 4203 6273 4212 6307
rect 4160 6264 4212 6273
rect 4620 6307 4672 6316
rect 4620 6273 4629 6307
rect 4629 6273 4663 6307
rect 4663 6273 4672 6307
rect 4620 6264 4672 6273
rect 5816 6264 5868 6316
rect 6736 6264 6788 6316
rect 7380 6264 7432 6316
rect 8852 6264 8904 6316
rect 9312 6400 9364 6452
rect 9404 6332 9456 6384
rect 9864 6400 9916 6452
rect 11244 6443 11296 6452
rect 11244 6409 11253 6443
rect 11253 6409 11287 6443
rect 11287 6409 11296 6443
rect 11244 6400 11296 6409
rect 4252 6196 4304 6248
rect 1860 6060 1912 6112
rect 3700 6128 3752 6180
rect 7932 6196 7984 6248
rect 8392 6196 8444 6248
rect 9588 6307 9640 6316
rect 9588 6273 9597 6307
rect 9597 6273 9631 6307
rect 9631 6273 9640 6307
rect 9588 6264 9640 6273
rect 9680 6293 9732 6316
rect 9680 6264 9689 6293
rect 9689 6264 9723 6293
rect 9723 6264 9732 6293
rect 10232 6332 10284 6384
rect 10508 6332 10560 6384
rect 10784 6332 10836 6384
rect 9312 6196 9364 6248
rect 10048 6307 10100 6316
rect 10048 6273 10057 6307
rect 10057 6273 10091 6307
rect 10091 6273 10100 6307
rect 10048 6264 10100 6273
rect 10692 6264 10744 6316
rect 11060 6307 11112 6316
rect 11060 6273 11069 6307
rect 11069 6273 11103 6307
rect 11103 6273 11112 6307
rect 11060 6264 11112 6273
rect 13176 6332 13228 6384
rect 10508 6196 10560 6248
rect 11796 6239 11848 6248
rect 11796 6205 11805 6239
rect 11805 6205 11839 6239
rect 11839 6205 11848 6239
rect 11796 6196 11848 6205
rect 8668 6128 8720 6180
rect 3608 6060 3660 6112
rect 3976 6060 4028 6112
rect 8484 6103 8536 6112
rect 8484 6069 8493 6103
rect 8493 6069 8527 6103
rect 8527 6069 8536 6103
rect 8484 6060 8536 6069
rect 9588 6060 9640 6112
rect 10600 6103 10652 6112
rect 10600 6069 10609 6103
rect 10609 6069 10643 6103
rect 10643 6069 10652 6103
rect 10600 6060 10652 6069
rect 10784 6103 10836 6112
rect 10784 6069 10793 6103
rect 10793 6069 10827 6103
rect 10827 6069 10836 6103
rect 10784 6060 10836 6069
rect 2525 5958 2577 6010
rect 2589 5958 2641 6010
rect 2653 5958 2705 6010
rect 2717 5958 2769 6010
rect 2781 5958 2833 6010
rect 5676 5958 5728 6010
rect 5740 5958 5792 6010
rect 5804 5958 5856 6010
rect 5868 5958 5920 6010
rect 5932 5958 5984 6010
rect 8827 5958 8879 6010
rect 8891 5958 8943 6010
rect 8955 5958 9007 6010
rect 9019 5958 9071 6010
rect 9083 5958 9135 6010
rect 11978 5958 12030 6010
rect 12042 5958 12094 6010
rect 12106 5958 12158 6010
rect 12170 5958 12222 6010
rect 12234 5958 12286 6010
rect 3516 5856 3568 5908
rect 4896 5856 4948 5908
rect 6184 5856 6236 5908
rect 10416 5899 10468 5908
rect 10416 5865 10425 5899
rect 10425 5865 10459 5899
rect 10459 5865 10468 5899
rect 10416 5856 10468 5865
rect 11796 5856 11848 5908
rect 4068 5788 4120 5840
rect 1768 5720 1820 5772
rect 2964 5720 3016 5772
rect 3424 5720 3476 5772
rect 2872 5652 2924 5704
rect 3700 5652 3752 5704
rect 3976 5695 4028 5704
rect 3976 5661 3985 5695
rect 3985 5661 4019 5695
rect 4019 5661 4028 5695
rect 3976 5652 4028 5661
rect 6828 5652 6880 5704
rect 10784 5652 10836 5704
rect 1768 5627 1820 5636
rect 1768 5593 1777 5627
rect 1777 5593 1811 5627
rect 1811 5593 1820 5627
rect 1768 5584 1820 5593
rect 4252 5584 4304 5636
rect 3185 5414 3237 5466
rect 3249 5414 3301 5466
rect 3313 5414 3365 5466
rect 3377 5414 3429 5466
rect 3441 5414 3493 5466
rect 6336 5414 6388 5466
rect 6400 5414 6452 5466
rect 6464 5414 6516 5466
rect 6528 5414 6580 5466
rect 6592 5414 6644 5466
rect 9487 5414 9539 5466
rect 9551 5414 9603 5466
rect 9615 5414 9667 5466
rect 9679 5414 9731 5466
rect 9743 5414 9795 5466
rect 12638 5414 12690 5466
rect 12702 5414 12754 5466
rect 12766 5414 12818 5466
rect 12830 5414 12882 5466
rect 12894 5414 12946 5466
rect 1768 5312 1820 5364
rect 3056 5312 3108 5364
rect 2872 5244 2924 5296
rect 4896 5287 4948 5296
rect 4896 5253 4905 5287
rect 4905 5253 4939 5287
rect 4939 5253 4948 5287
rect 4896 5244 4948 5253
rect 2136 5176 2188 5228
rect 3608 5176 3660 5228
rect 5540 5151 5592 5160
rect 5540 5117 5549 5151
rect 5549 5117 5583 5151
rect 5583 5117 5592 5151
rect 5540 5108 5592 5117
rect 6092 5040 6144 5092
rect 6000 5015 6052 5024
rect 6000 4981 6009 5015
rect 6009 4981 6043 5015
rect 6043 4981 6052 5015
rect 6000 4972 6052 4981
rect 9680 4972 9732 5024
rect 10784 4972 10836 5024
rect 2525 4870 2577 4922
rect 2589 4870 2641 4922
rect 2653 4870 2705 4922
rect 2717 4870 2769 4922
rect 2781 4870 2833 4922
rect 5676 4870 5728 4922
rect 5740 4870 5792 4922
rect 5804 4870 5856 4922
rect 5868 4870 5920 4922
rect 5932 4870 5984 4922
rect 8827 4870 8879 4922
rect 8891 4870 8943 4922
rect 8955 4870 9007 4922
rect 9019 4870 9071 4922
rect 9083 4870 9135 4922
rect 11978 4870 12030 4922
rect 12042 4870 12094 4922
rect 12106 4870 12158 4922
rect 12170 4870 12222 4922
rect 12234 4870 12286 4922
rect 3976 4768 4028 4820
rect 4804 4811 4856 4820
rect 4804 4777 4813 4811
rect 4813 4777 4847 4811
rect 4847 4777 4856 4811
rect 4804 4768 4856 4777
rect 3608 4700 3660 4752
rect 6828 4700 6880 4752
rect 4068 4632 4120 4684
rect 4896 4632 4948 4684
rect 5448 4675 5500 4684
rect 5448 4641 5457 4675
rect 5457 4641 5491 4675
rect 5491 4641 5500 4675
rect 5448 4632 5500 4641
rect 4344 4607 4396 4616
rect 4344 4573 4353 4607
rect 4353 4573 4387 4607
rect 4387 4573 4396 4607
rect 4344 4564 4396 4573
rect 4804 4564 4856 4616
rect 7932 4768 7984 4820
rect 8576 4632 8628 4684
rect 9956 4632 10008 4684
rect 10324 4675 10376 4684
rect 10324 4641 10333 4675
rect 10333 4641 10367 4675
rect 10367 4641 10376 4675
rect 10324 4632 10376 4641
rect 10968 4632 11020 4684
rect 9220 4564 9272 4616
rect 9312 4564 9364 4616
rect 9680 4607 9732 4616
rect 9680 4573 9689 4607
rect 9689 4573 9723 4607
rect 9723 4573 9732 4607
rect 9680 4564 9732 4573
rect 10048 4607 10100 4616
rect 10048 4573 10057 4607
rect 10057 4573 10091 4607
rect 10091 4573 10100 4607
rect 10048 4564 10100 4573
rect 12992 4564 13044 4616
rect 13176 4564 13228 4616
rect 4160 4471 4212 4480
rect 4160 4437 4169 4471
rect 4169 4437 4203 4471
rect 4203 4437 4212 4471
rect 4160 4428 4212 4437
rect 4620 4471 4672 4480
rect 4620 4437 4629 4471
rect 4629 4437 4663 4471
rect 4663 4437 4672 4471
rect 4620 4428 4672 4437
rect 4896 4428 4948 4480
rect 5632 4496 5684 4548
rect 5724 4539 5776 4548
rect 5724 4505 5733 4539
rect 5733 4505 5767 4539
rect 5767 4505 5776 4539
rect 5724 4496 5776 4505
rect 8300 4496 8352 4548
rect 10140 4496 10192 4548
rect 6092 4428 6144 4480
rect 8668 4428 8720 4480
rect 9128 4471 9180 4480
rect 9128 4437 9137 4471
rect 9137 4437 9171 4471
rect 9171 4437 9180 4471
rect 9128 4428 9180 4437
rect 9312 4428 9364 4480
rect 10784 4428 10836 4480
rect 12440 4428 12492 4480
rect 13084 4428 13136 4480
rect 13268 4471 13320 4480
rect 13268 4437 13277 4471
rect 13277 4437 13311 4471
rect 13311 4437 13320 4471
rect 13268 4428 13320 4437
rect 3185 4326 3237 4378
rect 3249 4326 3301 4378
rect 3313 4326 3365 4378
rect 3377 4326 3429 4378
rect 3441 4326 3493 4378
rect 6336 4326 6388 4378
rect 6400 4326 6452 4378
rect 6464 4326 6516 4378
rect 6528 4326 6580 4378
rect 6592 4326 6644 4378
rect 9487 4326 9539 4378
rect 9551 4326 9603 4378
rect 9615 4326 9667 4378
rect 9679 4326 9731 4378
rect 9743 4326 9795 4378
rect 12638 4326 12690 4378
rect 12702 4326 12754 4378
rect 12766 4326 12818 4378
rect 12830 4326 12882 4378
rect 12894 4326 12946 4378
rect 4344 4224 4396 4276
rect 5172 4224 5224 4276
rect 5540 4224 5592 4276
rect 5724 4224 5776 4276
rect 9956 4224 10008 4276
rect 10692 4224 10744 4276
rect 10968 4267 11020 4276
rect 10968 4233 10977 4267
rect 10977 4233 11011 4267
rect 11011 4233 11020 4267
rect 10968 4224 11020 4233
rect 5264 4131 5316 4140
rect 5264 4097 5273 4131
rect 5273 4097 5307 4131
rect 5307 4097 5316 4131
rect 5264 4088 5316 4097
rect 4252 3952 4304 4004
rect 5172 4020 5224 4072
rect 6000 4131 6052 4140
rect 6000 4097 6009 4131
rect 6009 4097 6043 4131
rect 6043 4097 6052 4131
rect 6000 4088 6052 4097
rect 6184 4156 6236 4208
rect 10324 4156 10376 4208
rect 10416 4156 10468 4208
rect 6828 4131 6880 4140
rect 6828 4097 6837 4131
rect 6837 4097 6871 4131
rect 6871 4097 6880 4131
rect 6828 4088 6880 4097
rect 3976 3884 4028 3936
rect 4988 3952 5040 4004
rect 5448 4020 5500 4072
rect 8392 4088 8444 4140
rect 9772 4131 9824 4140
rect 9772 4097 9781 4131
rect 9781 4097 9815 4131
rect 9815 4097 9824 4131
rect 9772 4088 9824 4097
rect 7656 4020 7708 4072
rect 9128 4020 9180 4072
rect 10140 4063 10192 4072
rect 10140 4029 10149 4063
rect 10149 4029 10183 4063
rect 10183 4029 10192 4063
rect 10140 4020 10192 4029
rect 10784 4088 10836 4140
rect 11152 4088 11204 4140
rect 12992 4131 13044 4140
rect 12992 4097 13001 4131
rect 13001 4097 13035 4131
rect 13035 4097 13044 4131
rect 12992 4088 13044 4097
rect 13084 4131 13136 4140
rect 13084 4097 13093 4131
rect 13093 4097 13127 4131
rect 13127 4097 13136 4131
rect 13084 4088 13136 4097
rect 5632 3952 5684 4004
rect 6000 3884 6052 3936
rect 6736 3952 6788 4004
rect 12532 3952 12584 4004
rect 13176 4020 13228 4072
rect 8300 3884 8352 3936
rect 9404 3884 9456 3936
rect 9956 3884 10008 3936
rect 11152 3927 11204 3936
rect 11152 3893 11161 3927
rect 11161 3893 11195 3927
rect 11195 3893 11204 3927
rect 11152 3884 11204 3893
rect 11520 3927 11572 3936
rect 11520 3893 11529 3927
rect 11529 3893 11563 3927
rect 11563 3893 11572 3927
rect 11520 3884 11572 3893
rect 2525 3782 2577 3834
rect 2589 3782 2641 3834
rect 2653 3782 2705 3834
rect 2717 3782 2769 3834
rect 2781 3782 2833 3834
rect 5676 3782 5728 3834
rect 5740 3782 5792 3834
rect 5804 3782 5856 3834
rect 5868 3782 5920 3834
rect 5932 3782 5984 3834
rect 8827 3782 8879 3834
rect 8891 3782 8943 3834
rect 8955 3782 9007 3834
rect 9019 3782 9071 3834
rect 9083 3782 9135 3834
rect 11978 3782 12030 3834
rect 12042 3782 12094 3834
rect 12106 3782 12158 3834
rect 12170 3782 12222 3834
rect 12234 3782 12286 3834
rect 848 3612 900 3664
rect 4620 3680 4672 3732
rect 5264 3680 5316 3732
rect 7656 3723 7708 3732
rect 7656 3689 7665 3723
rect 7665 3689 7699 3723
rect 7699 3689 7708 3723
rect 7656 3680 7708 3689
rect 10692 3723 10744 3732
rect 10692 3689 10701 3723
rect 10701 3689 10735 3723
rect 10735 3689 10744 3723
rect 10692 3680 10744 3689
rect 12532 3723 12584 3732
rect 12532 3689 12541 3723
rect 12541 3689 12575 3723
rect 12575 3689 12584 3723
rect 12532 3680 12584 3689
rect 3516 3544 3568 3596
rect 4068 3544 4120 3596
rect 5540 3544 5592 3596
rect 8484 3587 8536 3596
rect 8484 3553 8493 3587
rect 8493 3553 8527 3587
rect 8527 3553 8536 3587
rect 8484 3544 8536 3553
rect 9772 3544 9824 3596
rect 11520 3544 11572 3596
rect 3608 3476 3660 3528
rect 5816 3476 5868 3528
rect 7932 3519 7984 3528
rect 7932 3485 7941 3519
rect 7941 3485 7975 3519
rect 7975 3485 7984 3519
rect 7932 3476 7984 3485
rect 8576 3476 8628 3528
rect 13360 3519 13412 3528
rect 13360 3485 13369 3519
rect 13369 3485 13403 3519
rect 13403 3485 13412 3519
rect 13360 3476 13412 3485
rect 4068 3451 4120 3460
rect 4068 3417 4077 3451
rect 4077 3417 4111 3451
rect 4111 3417 4120 3451
rect 4068 3408 4120 3417
rect 3056 3340 3108 3392
rect 6920 3408 6972 3460
rect 12440 3408 12492 3460
rect 3185 3238 3237 3290
rect 3249 3238 3301 3290
rect 3313 3238 3365 3290
rect 3377 3238 3429 3290
rect 3441 3238 3493 3290
rect 6336 3238 6388 3290
rect 6400 3238 6452 3290
rect 6464 3238 6516 3290
rect 6528 3238 6580 3290
rect 6592 3238 6644 3290
rect 9487 3238 9539 3290
rect 9551 3238 9603 3290
rect 9615 3238 9667 3290
rect 9679 3238 9731 3290
rect 9743 3238 9795 3290
rect 12638 3238 12690 3290
rect 12702 3238 12754 3290
rect 12766 3238 12818 3290
rect 12830 3238 12882 3290
rect 12894 3238 12946 3290
rect 4896 3136 4948 3188
rect 5172 3136 5224 3188
rect 6092 3136 6144 3188
rect 6184 3136 6236 3188
rect 6920 3136 6972 3188
rect 8392 3136 8444 3188
rect 8668 3179 8720 3188
rect 8668 3145 8693 3179
rect 8693 3145 8720 3179
rect 8668 3136 8720 3145
rect 9220 3136 9272 3188
rect 9404 3136 9456 3188
rect 10048 3136 10100 3188
rect 3516 3068 3568 3120
rect 4160 3068 4212 3120
rect 848 2932 900 2984
rect 3056 2932 3108 2984
rect 4988 2932 5040 2984
rect 5448 3043 5500 3052
rect 5448 3009 5457 3043
rect 5457 3009 5491 3043
rect 5491 3009 5500 3043
rect 8484 3111 8536 3120
rect 8484 3077 8493 3111
rect 8493 3077 8527 3111
rect 8527 3077 8536 3111
rect 8484 3068 8536 3077
rect 5448 3000 5500 3009
rect 6828 3000 6880 3052
rect 7932 3000 7984 3052
rect 8576 3000 8628 3052
rect 11152 3000 11204 3052
rect 10232 2975 10284 2984
rect 10232 2941 10241 2975
rect 10241 2941 10275 2975
rect 10275 2941 10284 2975
rect 10232 2932 10284 2941
rect 10692 2932 10744 2984
rect 13360 2975 13412 2984
rect 13360 2941 13369 2975
rect 13369 2941 13403 2975
rect 13403 2941 13412 2975
rect 13360 2932 13412 2941
rect 9404 2864 9456 2916
rect 9312 2839 9364 2848
rect 9312 2805 9321 2839
rect 9321 2805 9355 2839
rect 9355 2805 9364 2839
rect 9312 2796 9364 2805
rect 2525 2694 2577 2746
rect 2589 2694 2641 2746
rect 2653 2694 2705 2746
rect 2717 2694 2769 2746
rect 2781 2694 2833 2746
rect 5676 2694 5728 2746
rect 5740 2694 5792 2746
rect 5804 2694 5856 2746
rect 5868 2694 5920 2746
rect 5932 2694 5984 2746
rect 8827 2694 8879 2746
rect 8891 2694 8943 2746
rect 8955 2694 9007 2746
rect 9019 2694 9071 2746
rect 9083 2694 9135 2746
rect 11978 2694 12030 2746
rect 12042 2694 12094 2746
rect 12106 2694 12158 2746
rect 12170 2694 12222 2746
rect 12234 2694 12286 2746
rect 4160 2635 4212 2644
rect 4160 2601 4169 2635
rect 4169 2601 4203 2635
rect 4203 2601 4212 2635
rect 4160 2592 4212 2601
rect 7380 2635 7432 2644
rect 7380 2601 7389 2635
rect 7389 2601 7423 2635
rect 7423 2601 7432 2635
rect 7380 2592 7432 2601
rect 3608 2388 3660 2440
rect 7104 2388 7156 2440
rect 10140 2456 10192 2508
rect 10232 2388 10284 2440
rect 10784 2388 10836 2440
rect 9036 2252 9088 2304
rect 9864 2295 9916 2304
rect 9864 2261 9873 2295
rect 9873 2261 9907 2295
rect 9907 2261 9916 2295
rect 9864 2252 9916 2261
rect 10324 2252 10376 2304
rect 3185 2150 3237 2202
rect 3249 2150 3301 2202
rect 3313 2150 3365 2202
rect 3377 2150 3429 2202
rect 3441 2150 3493 2202
rect 6336 2150 6388 2202
rect 6400 2150 6452 2202
rect 6464 2150 6516 2202
rect 6528 2150 6580 2202
rect 6592 2150 6644 2202
rect 9487 2150 9539 2202
rect 9551 2150 9603 2202
rect 9615 2150 9667 2202
rect 9679 2150 9731 2202
rect 9743 2150 9795 2202
rect 12638 2150 12690 2202
rect 12702 2150 12754 2202
rect 12766 2150 12818 2202
rect 12830 2150 12882 2202
rect 12894 2150 12946 2202
<< metal2 >>
rect 2525 14716 2833 14725
rect 2525 14714 2531 14716
rect 2587 14714 2611 14716
rect 2667 14714 2691 14716
rect 2747 14714 2771 14716
rect 2827 14714 2833 14716
rect 2587 14662 2589 14714
rect 2769 14662 2771 14714
rect 2525 14660 2531 14662
rect 2587 14660 2611 14662
rect 2667 14660 2691 14662
rect 2747 14660 2771 14662
rect 2827 14660 2833 14662
rect 2525 14651 2833 14660
rect 5676 14716 5984 14725
rect 5676 14714 5682 14716
rect 5738 14714 5762 14716
rect 5818 14714 5842 14716
rect 5898 14714 5922 14716
rect 5978 14714 5984 14716
rect 5738 14662 5740 14714
rect 5920 14662 5922 14714
rect 5676 14660 5682 14662
rect 5738 14660 5762 14662
rect 5818 14660 5842 14662
rect 5898 14660 5922 14662
rect 5978 14660 5984 14662
rect 5676 14651 5984 14660
rect 8827 14716 9135 14725
rect 8827 14714 8833 14716
rect 8889 14714 8913 14716
rect 8969 14714 8993 14716
rect 9049 14714 9073 14716
rect 9129 14714 9135 14716
rect 8889 14662 8891 14714
rect 9071 14662 9073 14714
rect 8827 14660 8833 14662
rect 8889 14660 8913 14662
rect 8969 14660 8993 14662
rect 9049 14660 9073 14662
rect 9129 14660 9135 14662
rect 8827 14651 9135 14660
rect 11978 14716 12286 14725
rect 11978 14714 11984 14716
rect 12040 14714 12064 14716
rect 12120 14714 12144 14716
rect 12200 14714 12224 14716
rect 12280 14714 12286 14716
rect 12040 14662 12042 14714
rect 12222 14662 12224 14714
rect 11978 14660 11984 14662
rect 12040 14660 12064 14662
rect 12120 14660 12144 14662
rect 12200 14660 12224 14662
rect 12280 14660 12286 14662
rect 11978 14651 12286 14660
rect 3185 14172 3493 14181
rect 3185 14170 3191 14172
rect 3247 14170 3271 14172
rect 3327 14170 3351 14172
rect 3407 14170 3431 14172
rect 3487 14170 3493 14172
rect 3247 14118 3249 14170
rect 3429 14118 3431 14170
rect 3185 14116 3191 14118
rect 3247 14116 3271 14118
rect 3327 14116 3351 14118
rect 3407 14116 3431 14118
rect 3487 14116 3493 14118
rect 3185 14107 3493 14116
rect 6336 14172 6644 14181
rect 6336 14170 6342 14172
rect 6398 14170 6422 14172
rect 6478 14170 6502 14172
rect 6558 14170 6582 14172
rect 6638 14170 6644 14172
rect 6398 14118 6400 14170
rect 6580 14118 6582 14170
rect 6336 14116 6342 14118
rect 6398 14116 6422 14118
rect 6478 14116 6502 14118
rect 6558 14116 6582 14118
rect 6638 14116 6644 14118
rect 6336 14107 6644 14116
rect 9487 14172 9795 14181
rect 9487 14170 9493 14172
rect 9549 14170 9573 14172
rect 9629 14170 9653 14172
rect 9709 14170 9733 14172
rect 9789 14170 9795 14172
rect 9549 14118 9551 14170
rect 9731 14118 9733 14170
rect 9487 14116 9493 14118
rect 9549 14116 9573 14118
rect 9629 14116 9653 14118
rect 9709 14116 9733 14118
rect 9789 14116 9795 14118
rect 9487 14107 9795 14116
rect 12638 14172 12946 14181
rect 12638 14170 12644 14172
rect 12700 14170 12724 14172
rect 12780 14170 12804 14172
rect 12860 14170 12884 14172
rect 12940 14170 12946 14172
rect 12700 14118 12702 14170
rect 12882 14118 12884 14170
rect 12638 14116 12644 14118
rect 12700 14116 12724 14118
rect 12780 14116 12804 14118
rect 12860 14116 12884 14118
rect 12940 14116 12946 14118
rect 12638 14107 12946 14116
rect 9588 14000 9640 14006
rect 9588 13942 9640 13948
rect 6460 13932 6512 13938
rect 6460 13874 6512 13880
rect 6736 13932 6788 13938
rect 6736 13874 6788 13880
rect 1400 13864 1452 13870
rect 1400 13806 1452 13812
rect 5816 13864 5868 13870
rect 5868 13812 6040 13818
rect 5816 13806 6040 13812
rect 1412 13705 1440 13806
rect 5540 13796 5592 13802
rect 5828 13790 6040 13806
rect 5540 13738 5592 13744
rect 4620 13728 4672 13734
rect 1398 13696 1454 13705
rect 4620 13670 4672 13676
rect 5448 13728 5500 13734
rect 5448 13670 5500 13676
rect 1398 13631 1454 13640
rect 2525 13628 2833 13637
rect 2525 13626 2531 13628
rect 2587 13626 2611 13628
rect 2667 13626 2691 13628
rect 2747 13626 2771 13628
rect 2827 13626 2833 13628
rect 2587 13574 2589 13626
rect 2769 13574 2771 13626
rect 2525 13572 2531 13574
rect 2587 13572 2611 13574
rect 2667 13572 2691 13574
rect 2747 13572 2771 13574
rect 2827 13572 2833 13574
rect 2525 13563 2833 13572
rect 4160 13388 4212 13394
rect 4160 13330 4212 13336
rect 3700 13320 3752 13326
rect 3700 13262 3752 13268
rect 848 13184 900 13190
rect 846 13152 848 13161
rect 2872 13184 2924 13190
rect 900 13152 902 13161
rect 2872 13126 2924 13132
rect 3516 13184 3568 13190
rect 3516 13126 3568 13132
rect 846 13087 902 13096
rect 2884 12918 2912 13126
rect 3185 13084 3493 13093
rect 3185 13082 3191 13084
rect 3247 13082 3271 13084
rect 3327 13082 3351 13084
rect 3407 13082 3431 13084
rect 3487 13082 3493 13084
rect 3247 13030 3249 13082
rect 3429 13030 3431 13082
rect 3185 13028 3191 13030
rect 3247 13028 3271 13030
rect 3327 13028 3351 13030
rect 3407 13028 3431 13030
rect 3487 13028 3493 13030
rect 3185 13019 3493 13028
rect 3528 12918 3556 13126
rect 2872 12912 2924 12918
rect 2872 12854 2924 12860
rect 3516 12912 3568 12918
rect 3516 12854 3568 12860
rect 1676 12776 1728 12782
rect 1676 12718 1728 12724
rect 1688 11898 1716 12718
rect 2525 12540 2833 12549
rect 2525 12538 2531 12540
rect 2587 12538 2611 12540
rect 2667 12538 2691 12540
rect 2747 12538 2771 12540
rect 2827 12538 2833 12540
rect 2587 12486 2589 12538
rect 2769 12486 2771 12538
rect 2525 12484 2531 12486
rect 2587 12484 2611 12486
rect 2667 12484 2691 12486
rect 2747 12484 2771 12486
rect 2827 12484 2833 12486
rect 2525 12475 2833 12484
rect 3185 11996 3493 12005
rect 3185 11994 3191 11996
rect 3247 11994 3271 11996
rect 3327 11994 3351 11996
rect 3407 11994 3431 11996
rect 3487 11994 3493 11996
rect 3247 11942 3249 11994
rect 3429 11942 3431 11994
rect 3185 11940 3191 11942
rect 3247 11940 3271 11942
rect 3327 11940 3351 11942
rect 3407 11940 3431 11942
rect 3487 11940 3493 11942
rect 3185 11931 3493 11940
rect 1676 11892 1728 11898
rect 1676 11834 1728 11840
rect 1688 11694 1716 11834
rect 3712 11762 3740 13262
rect 4172 12782 4200 13330
rect 4632 13258 4660 13670
rect 4804 13524 4856 13530
rect 4804 13466 4856 13472
rect 4816 13326 4844 13466
rect 4804 13320 4856 13326
rect 4804 13262 4856 13268
rect 4528 13252 4580 13258
rect 4528 13194 4580 13200
rect 4620 13252 4672 13258
rect 4620 13194 4672 13200
rect 4344 13184 4396 13190
rect 4344 13126 4396 13132
rect 4160 12776 4212 12782
rect 4160 12718 4212 12724
rect 4172 12434 4200 12718
rect 4356 12442 4384 13126
rect 4344 12436 4396 12442
rect 4172 12406 4292 12434
rect 4160 12096 4212 12102
rect 4160 12038 4212 12044
rect 3700 11756 3752 11762
rect 3700 11698 3752 11704
rect 1676 11688 1728 11694
rect 1676 11630 1728 11636
rect 1952 11688 2004 11694
rect 1952 11630 2004 11636
rect 1492 10668 1544 10674
rect 1492 10610 1544 10616
rect 1504 10266 1532 10610
rect 1688 10606 1716 11630
rect 1964 11354 1992 11630
rect 3712 11626 3740 11698
rect 3700 11620 3752 11626
rect 3700 11562 3752 11568
rect 2525 11452 2833 11461
rect 2525 11450 2531 11452
rect 2587 11450 2611 11452
rect 2667 11450 2691 11452
rect 2747 11450 2771 11452
rect 2827 11450 2833 11452
rect 2587 11398 2589 11450
rect 2769 11398 2771 11450
rect 2525 11396 2531 11398
rect 2587 11396 2611 11398
rect 2667 11396 2691 11398
rect 2747 11396 2771 11398
rect 2827 11396 2833 11398
rect 2525 11387 2833 11396
rect 1952 11348 2004 11354
rect 1952 11290 2004 11296
rect 2964 11144 3016 11150
rect 2964 11086 3016 11092
rect 2412 11008 2464 11014
rect 2412 10950 2464 10956
rect 2872 11008 2924 11014
rect 2872 10950 2924 10956
rect 1676 10600 1728 10606
rect 1676 10542 1728 10548
rect 1492 10260 1544 10266
rect 1492 10202 1544 10208
rect 1688 8498 1716 10542
rect 2424 10062 2452 10950
rect 2525 10364 2833 10373
rect 2525 10362 2531 10364
rect 2587 10362 2611 10364
rect 2667 10362 2691 10364
rect 2747 10362 2771 10364
rect 2827 10362 2833 10364
rect 2587 10310 2589 10362
rect 2769 10310 2771 10362
rect 2525 10308 2531 10310
rect 2587 10308 2611 10310
rect 2667 10308 2691 10310
rect 2747 10308 2771 10310
rect 2827 10308 2833 10310
rect 2525 10299 2833 10308
rect 2412 10056 2464 10062
rect 2412 9998 2464 10004
rect 2884 9926 2912 10950
rect 2976 10266 3004 11086
rect 3185 10908 3493 10917
rect 3185 10906 3191 10908
rect 3247 10906 3271 10908
rect 3327 10906 3351 10908
rect 3407 10906 3431 10908
rect 3487 10906 3493 10908
rect 3247 10854 3249 10906
rect 3429 10854 3431 10906
rect 3185 10852 3191 10854
rect 3247 10852 3271 10854
rect 3327 10852 3351 10854
rect 3407 10852 3431 10854
rect 3487 10852 3493 10854
rect 3185 10843 3493 10852
rect 3056 10736 3108 10742
rect 3056 10678 3108 10684
rect 2964 10260 3016 10266
rect 2964 10202 3016 10208
rect 2872 9920 2924 9926
rect 2872 9862 2924 9868
rect 2964 9920 3016 9926
rect 2964 9862 3016 9868
rect 2872 9512 2924 9518
rect 2872 9454 2924 9460
rect 2525 9276 2833 9285
rect 2525 9274 2531 9276
rect 2587 9274 2611 9276
rect 2667 9274 2691 9276
rect 2747 9274 2771 9276
rect 2827 9274 2833 9276
rect 2587 9222 2589 9274
rect 2769 9222 2771 9274
rect 2525 9220 2531 9222
rect 2587 9220 2611 9222
rect 2667 9220 2691 9222
rect 2747 9220 2771 9222
rect 2827 9220 2833 9222
rect 2525 9211 2833 9220
rect 1952 8832 2004 8838
rect 1952 8774 2004 8780
rect 1964 8566 1992 8774
rect 1952 8560 2004 8566
rect 1952 8502 2004 8508
rect 1676 8492 1728 8498
rect 1676 8434 1728 8440
rect 2525 8188 2833 8197
rect 2525 8186 2531 8188
rect 2587 8186 2611 8188
rect 2667 8186 2691 8188
rect 2747 8186 2771 8188
rect 2827 8186 2833 8188
rect 2587 8134 2589 8186
rect 2769 8134 2771 8186
rect 2525 8132 2531 8134
rect 2587 8132 2611 8134
rect 2667 8132 2691 8134
rect 2747 8132 2771 8134
rect 2827 8132 2833 8134
rect 2525 8123 2833 8132
rect 2884 7886 2912 9454
rect 2976 8906 3004 9862
rect 3068 9654 3096 10678
rect 3424 10464 3476 10470
rect 3424 10406 3476 10412
rect 3332 10260 3384 10266
rect 3332 10202 3384 10208
rect 3344 10062 3372 10202
rect 3436 10062 3464 10406
rect 3332 10056 3384 10062
rect 3332 9998 3384 10004
rect 3424 10056 3476 10062
rect 3424 9998 3476 10004
rect 3185 9820 3493 9829
rect 3185 9818 3191 9820
rect 3247 9818 3271 9820
rect 3327 9818 3351 9820
rect 3407 9818 3431 9820
rect 3487 9818 3493 9820
rect 3247 9766 3249 9818
rect 3429 9766 3431 9818
rect 3185 9764 3191 9766
rect 3247 9764 3271 9766
rect 3327 9764 3351 9766
rect 3407 9764 3431 9766
rect 3487 9764 3493 9766
rect 3185 9755 3493 9764
rect 3712 9654 3740 11562
rect 3792 11552 3844 11558
rect 3792 11494 3844 11500
rect 3804 10742 3832 11494
rect 4172 11234 4200 12038
rect 4264 11898 4292 12406
rect 4344 12378 4396 12384
rect 4540 12102 4568 13194
rect 4816 12986 4844 13262
rect 5080 13184 5132 13190
rect 5080 13126 5132 13132
rect 4804 12980 4856 12986
rect 4804 12922 4856 12928
rect 4712 12776 4764 12782
rect 4712 12718 4764 12724
rect 4724 12442 4752 12718
rect 4712 12436 4764 12442
rect 4712 12378 4764 12384
rect 4620 12368 4672 12374
rect 4620 12310 4672 12316
rect 4528 12096 4580 12102
rect 4528 12038 4580 12044
rect 4252 11892 4304 11898
rect 4252 11834 4304 11840
rect 4264 11558 4292 11834
rect 4252 11552 4304 11558
rect 4252 11494 4304 11500
rect 4080 11206 4200 11234
rect 3792 10736 3844 10742
rect 3792 10678 3844 10684
rect 3804 10266 3832 10678
rect 3792 10260 3844 10266
rect 3792 10202 3844 10208
rect 4080 9926 4108 11206
rect 4160 11144 4212 11150
rect 4160 11086 4212 11092
rect 4172 10810 4200 11086
rect 4264 11082 4292 11494
rect 4632 11150 4660 12310
rect 5092 12238 5120 13126
rect 5460 12374 5488 13670
rect 5552 13190 5580 13738
rect 5676 13628 5984 13637
rect 5676 13626 5682 13628
rect 5738 13626 5762 13628
rect 5818 13626 5842 13628
rect 5898 13626 5922 13628
rect 5978 13626 5984 13628
rect 5738 13574 5740 13626
rect 5920 13574 5922 13626
rect 5676 13572 5682 13574
rect 5738 13572 5762 13574
rect 5818 13572 5842 13574
rect 5898 13572 5922 13574
rect 5978 13572 5984 13574
rect 5676 13563 5984 13572
rect 6012 13530 6040 13790
rect 6184 13728 6236 13734
rect 6184 13670 6236 13676
rect 6368 13728 6420 13734
rect 6368 13670 6420 13676
rect 6000 13524 6052 13530
rect 6000 13466 6052 13472
rect 5540 13184 5592 13190
rect 5540 13126 5592 13132
rect 5552 12986 5580 13126
rect 5540 12980 5592 12986
rect 5540 12922 5592 12928
rect 6012 12850 6040 13466
rect 6092 12980 6144 12986
rect 6092 12922 6144 12928
rect 6000 12844 6052 12850
rect 6000 12786 6052 12792
rect 5676 12540 5984 12549
rect 5676 12538 5682 12540
rect 5738 12538 5762 12540
rect 5818 12538 5842 12540
rect 5898 12538 5922 12540
rect 5978 12538 5984 12540
rect 5738 12486 5740 12538
rect 5920 12486 5922 12538
rect 5676 12484 5682 12486
rect 5738 12484 5762 12486
rect 5818 12484 5842 12486
rect 5898 12484 5922 12486
rect 5978 12484 5984 12486
rect 5676 12475 5984 12484
rect 6012 12434 6040 12786
rect 6104 12646 6132 12922
rect 6092 12640 6144 12646
rect 6092 12582 6144 12588
rect 5920 12406 6040 12434
rect 5448 12368 5500 12374
rect 5448 12310 5500 12316
rect 5080 12232 5132 12238
rect 5080 12174 5132 12180
rect 5172 12232 5224 12238
rect 5172 12174 5224 12180
rect 5448 12232 5500 12238
rect 5448 12174 5500 12180
rect 5184 11830 5212 12174
rect 5172 11824 5224 11830
rect 5172 11766 5224 11772
rect 4896 11552 4948 11558
rect 4896 11494 4948 11500
rect 4908 11150 4936 11494
rect 5184 11354 5212 11766
rect 5172 11348 5224 11354
rect 5172 11290 5224 11296
rect 4620 11144 4672 11150
rect 4896 11144 4948 11150
rect 4672 11104 4752 11132
rect 4620 11086 4672 11092
rect 4252 11076 4304 11082
rect 4252 11018 4304 11024
rect 4528 11008 4580 11014
rect 4528 10950 4580 10956
rect 4620 11008 4672 11014
rect 4620 10950 4672 10956
rect 4160 10804 4212 10810
rect 4160 10746 4212 10752
rect 4160 10668 4212 10674
rect 4160 10610 4212 10616
rect 4172 9926 4200 10610
rect 4540 10606 4568 10950
rect 4528 10600 4580 10606
rect 4528 10542 4580 10548
rect 4436 10532 4488 10538
rect 4436 10474 4488 10480
rect 4344 10464 4396 10470
rect 4344 10406 4396 10412
rect 4252 10124 4304 10130
rect 4252 10066 4304 10072
rect 4068 9920 4120 9926
rect 4068 9862 4120 9868
rect 4160 9920 4212 9926
rect 4160 9862 4212 9868
rect 3056 9648 3108 9654
rect 3056 9590 3108 9596
rect 3700 9648 3752 9654
rect 3700 9590 3752 9596
rect 4172 9586 4200 9862
rect 4264 9654 4292 10066
rect 4356 10062 4384 10406
rect 4448 10062 4476 10474
rect 4344 10056 4396 10062
rect 4344 9998 4396 10004
rect 4436 10056 4488 10062
rect 4436 9998 4488 10004
rect 4252 9648 4304 9654
rect 4252 9590 4304 9596
rect 4160 9580 4212 9586
rect 4160 9522 4212 9528
rect 4344 9580 4396 9586
rect 4344 9522 4396 9528
rect 4436 9580 4488 9586
rect 4436 9522 4488 9528
rect 3884 9444 3936 9450
rect 3884 9386 3936 9392
rect 3148 9376 3200 9382
rect 3148 9318 3200 9324
rect 3160 9178 3188 9318
rect 3148 9172 3200 9178
rect 3148 9114 3200 9120
rect 3896 8906 3924 9386
rect 4172 9178 4200 9522
rect 4160 9172 4212 9178
rect 4160 9114 4212 9120
rect 4356 9110 4384 9522
rect 4344 9104 4396 9110
rect 4344 9046 4396 9052
rect 4448 8906 4476 9522
rect 4540 9518 4568 10542
rect 4632 9994 4660 10950
rect 4724 10538 4752 11104
rect 4896 11086 4948 11092
rect 5172 11144 5224 11150
rect 5172 11086 5224 11092
rect 4804 10600 4856 10606
rect 4804 10542 4856 10548
rect 4712 10532 4764 10538
rect 4712 10474 4764 10480
rect 4816 10282 4844 10542
rect 4724 10266 4844 10282
rect 4712 10260 4844 10266
rect 4764 10254 4844 10260
rect 4712 10202 4764 10208
rect 4620 9988 4672 9994
rect 4620 9930 4672 9936
rect 4528 9512 4580 9518
rect 4528 9454 4580 9460
rect 4632 9330 4660 9930
rect 4816 9382 4844 10254
rect 5184 10130 5212 11086
rect 5460 11014 5488 12174
rect 5920 12170 5948 12406
rect 6104 12306 6132 12582
rect 6196 12442 6224 13670
rect 6380 13394 6408 13670
rect 6472 13530 6500 13874
rect 6460 13524 6512 13530
rect 6460 13466 6512 13472
rect 6368 13388 6420 13394
rect 6368 13330 6420 13336
rect 6336 13084 6644 13093
rect 6336 13082 6342 13084
rect 6398 13082 6422 13084
rect 6478 13082 6502 13084
rect 6558 13082 6582 13084
rect 6638 13082 6644 13084
rect 6398 13030 6400 13082
rect 6580 13030 6582 13082
rect 6336 13028 6342 13030
rect 6398 13028 6422 13030
rect 6478 13028 6502 13030
rect 6558 13028 6582 13030
rect 6638 13028 6644 13030
rect 6336 13019 6644 13028
rect 6748 12442 6776 13874
rect 9496 13864 9548 13870
rect 9496 13806 9548 13812
rect 7932 13728 7984 13734
rect 7932 13670 7984 13676
rect 6828 13524 6880 13530
rect 6828 13466 6880 13472
rect 7840 13524 7892 13530
rect 7840 13466 7892 13472
rect 6840 12918 6868 13466
rect 7104 13320 7156 13326
rect 7104 13262 7156 13268
rect 6828 12912 6880 12918
rect 6828 12854 6880 12860
rect 7116 12850 7144 13262
rect 7196 13252 7248 13258
rect 7196 13194 7248 13200
rect 7104 12844 7156 12850
rect 7104 12786 7156 12792
rect 6828 12640 6880 12646
rect 6828 12582 6880 12588
rect 6920 12640 6972 12646
rect 6920 12582 6972 12588
rect 6184 12436 6236 12442
rect 6184 12378 6236 12384
rect 6736 12436 6788 12442
rect 6736 12378 6788 12384
rect 6092 12300 6144 12306
rect 6092 12242 6144 12248
rect 5908 12164 5960 12170
rect 5908 12106 5960 12112
rect 6184 12096 6236 12102
rect 6184 12038 6236 12044
rect 6196 11830 6224 12038
rect 6336 11996 6644 12005
rect 6336 11994 6342 11996
rect 6398 11994 6422 11996
rect 6478 11994 6502 11996
rect 6558 11994 6582 11996
rect 6638 11994 6644 11996
rect 6398 11942 6400 11994
rect 6580 11942 6582 11994
rect 6336 11940 6342 11942
rect 6398 11940 6422 11942
rect 6478 11940 6502 11942
rect 6558 11940 6582 11942
rect 6638 11940 6644 11942
rect 6336 11931 6644 11940
rect 6184 11824 6236 11830
rect 6184 11766 6236 11772
rect 6552 11756 6604 11762
rect 6552 11698 6604 11704
rect 5540 11688 5592 11694
rect 5540 11630 5592 11636
rect 5448 11008 5500 11014
rect 5448 10950 5500 10956
rect 5552 10810 5580 11630
rect 5676 11452 5984 11461
rect 5676 11450 5682 11452
rect 5738 11450 5762 11452
rect 5818 11450 5842 11452
rect 5898 11450 5922 11452
rect 5978 11450 5984 11452
rect 5738 11398 5740 11450
rect 5920 11398 5922 11450
rect 5676 11396 5682 11398
rect 5738 11396 5762 11398
rect 5818 11396 5842 11398
rect 5898 11396 5922 11398
rect 5978 11396 5984 11398
rect 5676 11387 5984 11396
rect 6564 11354 6592 11698
rect 5908 11348 5960 11354
rect 5908 11290 5960 11296
rect 6552 11348 6604 11354
rect 6552 11290 6604 11296
rect 5540 10804 5592 10810
rect 5540 10746 5592 10752
rect 5920 10742 5948 11290
rect 6336 10908 6644 10917
rect 6336 10906 6342 10908
rect 6398 10906 6422 10908
rect 6478 10906 6502 10908
rect 6558 10906 6582 10908
rect 6638 10906 6644 10908
rect 6398 10854 6400 10906
rect 6580 10854 6582 10906
rect 6336 10852 6342 10854
rect 6398 10852 6422 10854
rect 6478 10852 6502 10854
rect 6558 10852 6582 10854
rect 6638 10852 6644 10854
rect 6336 10843 6644 10852
rect 5908 10736 5960 10742
rect 6840 10690 6868 12582
rect 6932 12170 6960 12582
rect 6920 12164 6972 12170
rect 6920 12106 6972 12112
rect 7116 11762 7144 12786
rect 7208 12102 7236 13194
rect 7748 13184 7800 13190
rect 7748 13126 7800 13132
rect 7760 12850 7788 13126
rect 7852 12986 7880 13466
rect 7840 12980 7892 12986
rect 7840 12922 7892 12928
rect 7944 12866 7972 13670
rect 8827 13628 9135 13637
rect 8827 13626 8833 13628
rect 8889 13626 8913 13628
rect 8969 13626 8993 13628
rect 9049 13626 9073 13628
rect 9129 13626 9135 13628
rect 8889 13574 8891 13626
rect 9071 13574 9073 13626
rect 8827 13572 8833 13574
rect 8889 13572 8913 13574
rect 8969 13572 8993 13574
rect 9049 13572 9073 13574
rect 9129 13572 9135 13574
rect 8827 13563 9135 13572
rect 9508 13530 9536 13806
rect 9600 13530 9628 13942
rect 10232 13864 10284 13870
rect 10232 13806 10284 13812
rect 13360 13864 13412 13870
rect 13360 13806 13412 13812
rect 9496 13524 9548 13530
rect 9496 13466 9548 13472
rect 9588 13524 9640 13530
rect 9588 13466 9640 13472
rect 8392 13320 8444 13326
rect 8392 13262 8444 13268
rect 9128 13320 9180 13326
rect 9128 13262 9180 13268
rect 8208 13252 8260 13258
rect 8208 13194 8260 13200
rect 7944 12850 8064 12866
rect 7748 12844 7800 12850
rect 7748 12786 7800 12792
rect 7932 12844 8064 12850
rect 7984 12838 8064 12844
rect 7932 12786 7984 12792
rect 7932 12708 7984 12714
rect 7932 12650 7984 12656
rect 7944 12306 7972 12650
rect 8036 12646 8064 12838
rect 8024 12640 8076 12646
rect 8024 12582 8076 12588
rect 8220 12442 8248 13194
rect 8404 12986 8432 13262
rect 8484 13252 8536 13258
rect 8484 13194 8536 13200
rect 8496 12986 8524 13194
rect 8576 13184 8628 13190
rect 8576 13126 8628 13132
rect 8392 12980 8444 12986
rect 8392 12922 8444 12928
rect 8484 12980 8536 12986
rect 8484 12922 8536 12928
rect 8392 12640 8444 12646
rect 8392 12582 8444 12588
rect 8208 12436 8260 12442
rect 8208 12378 8260 12384
rect 7932 12300 7984 12306
rect 7932 12242 7984 12248
rect 7196 12096 7248 12102
rect 7196 12038 7248 12044
rect 7104 11756 7156 11762
rect 7104 11698 7156 11704
rect 6920 11552 6972 11558
rect 6920 11494 6972 11500
rect 6932 11150 6960 11494
rect 6920 11144 6972 11150
rect 6920 11086 6972 11092
rect 5908 10678 5960 10684
rect 5264 10668 5316 10674
rect 5264 10610 5316 10616
rect 5356 10668 5408 10674
rect 5356 10610 5408 10616
rect 5172 10124 5224 10130
rect 5172 10066 5224 10072
rect 5276 9722 5304 10610
rect 5368 10538 5396 10610
rect 5920 10606 5948 10678
rect 6748 10674 6868 10690
rect 6736 10668 6868 10674
rect 6788 10662 6868 10668
rect 6736 10610 6788 10616
rect 5908 10600 5960 10606
rect 5908 10542 5960 10548
rect 5356 10532 5408 10538
rect 5356 10474 5408 10480
rect 5368 9926 5396 10474
rect 5676 10364 5984 10373
rect 5676 10362 5682 10364
rect 5738 10362 5762 10364
rect 5818 10362 5842 10364
rect 5898 10362 5922 10364
rect 5978 10362 5984 10364
rect 5738 10310 5740 10362
rect 5920 10310 5922 10362
rect 5676 10308 5682 10310
rect 5738 10308 5762 10310
rect 5818 10308 5842 10310
rect 5898 10308 5922 10310
rect 5978 10308 5984 10310
rect 5676 10299 5984 10308
rect 5356 9920 5408 9926
rect 5356 9862 5408 9868
rect 5264 9716 5316 9722
rect 5264 9658 5316 9664
rect 5368 9654 5396 9862
rect 6336 9820 6644 9829
rect 6336 9818 6342 9820
rect 6398 9818 6422 9820
rect 6478 9818 6502 9820
rect 6558 9818 6582 9820
rect 6638 9818 6644 9820
rect 6398 9766 6400 9818
rect 6580 9766 6582 9818
rect 6336 9764 6342 9766
rect 6398 9764 6422 9766
rect 6478 9764 6502 9766
rect 6558 9764 6582 9766
rect 6638 9764 6644 9766
rect 6336 9755 6644 9764
rect 5356 9648 5408 9654
rect 5356 9590 5408 9596
rect 6550 9616 6606 9625
rect 6550 9551 6606 9560
rect 4540 9302 4660 9330
rect 4804 9376 4856 9382
rect 4804 9318 4856 9324
rect 5356 9376 5408 9382
rect 5356 9318 5408 9324
rect 2964 8900 3016 8906
rect 2964 8842 3016 8848
rect 3884 8900 3936 8906
rect 3884 8842 3936 8848
rect 4436 8900 4488 8906
rect 4436 8842 4488 8848
rect 2976 8650 3004 8842
rect 3516 8832 3568 8838
rect 3516 8774 3568 8780
rect 3185 8732 3493 8741
rect 3185 8730 3191 8732
rect 3247 8730 3271 8732
rect 3327 8730 3351 8732
rect 3407 8730 3431 8732
rect 3487 8730 3493 8732
rect 3247 8678 3249 8730
rect 3429 8678 3431 8730
rect 3185 8676 3191 8678
rect 3247 8676 3271 8678
rect 3327 8676 3351 8678
rect 3407 8676 3431 8678
rect 3487 8676 3493 8678
rect 3185 8667 3493 8676
rect 2976 8622 3096 8650
rect 3528 8634 3556 8774
rect 3896 8634 3924 8842
rect 2964 8560 3016 8566
rect 2964 8502 3016 8508
rect 2976 8090 3004 8502
rect 2964 8084 3016 8090
rect 2964 8026 3016 8032
rect 2872 7880 2924 7886
rect 2872 7822 2924 7828
rect 2320 7200 2372 7206
rect 2320 7142 2372 7148
rect 2332 7002 2360 7142
rect 2525 7100 2833 7109
rect 2525 7098 2531 7100
rect 2587 7098 2611 7100
rect 2667 7098 2691 7100
rect 2747 7098 2771 7100
rect 2827 7098 2833 7100
rect 2587 7046 2589 7098
rect 2769 7046 2771 7098
rect 2525 7044 2531 7046
rect 2587 7044 2611 7046
rect 2667 7044 2691 7046
rect 2747 7044 2771 7046
rect 2827 7044 2833 7046
rect 2525 7035 2833 7044
rect 2320 6996 2372 7002
rect 2320 6938 2372 6944
rect 2964 6996 3016 7002
rect 2964 6938 3016 6944
rect 2136 6928 2188 6934
rect 2136 6870 2188 6876
rect 1860 6792 1912 6798
rect 1860 6734 1912 6740
rect 1492 6724 1544 6730
rect 1492 6666 1544 6672
rect 1504 6322 1532 6666
rect 1492 6316 1544 6322
rect 1492 6258 1544 6264
rect 1768 6316 1820 6322
rect 1768 6258 1820 6264
rect 1780 5778 1808 6258
rect 1872 6118 1900 6734
rect 1860 6112 1912 6118
rect 1860 6054 1912 6060
rect 1768 5772 1820 5778
rect 1768 5714 1820 5720
rect 1768 5636 1820 5642
rect 1768 5578 1820 5584
rect 1780 5370 1808 5578
rect 1768 5364 1820 5370
rect 1768 5306 1820 5312
rect 2148 5234 2176 6870
rect 2516 6866 2728 6882
rect 2504 6860 2740 6866
rect 2556 6854 2688 6860
rect 2504 6802 2556 6808
rect 2688 6802 2740 6808
rect 2525 6012 2833 6021
rect 2525 6010 2531 6012
rect 2587 6010 2611 6012
rect 2667 6010 2691 6012
rect 2747 6010 2771 6012
rect 2827 6010 2833 6012
rect 2587 5958 2589 6010
rect 2769 5958 2771 6010
rect 2525 5956 2531 5958
rect 2587 5956 2611 5958
rect 2667 5956 2691 5958
rect 2747 5956 2771 5958
rect 2827 5956 2833 5958
rect 2525 5947 2833 5956
rect 2976 5778 3004 6938
rect 3068 6730 3096 8622
rect 3516 8628 3568 8634
rect 3516 8570 3568 8576
rect 3884 8628 3936 8634
rect 3884 8570 3936 8576
rect 4344 8492 4396 8498
rect 4344 8434 4396 8440
rect 4356 8022 4384 8434
rect 4344 8016 4396 8022
rect 4344 7958 4396 7964
rect 4436 7812 4488 7818
rect 4436 7754 4488 7760
rect 3185 7644 3493 7653
rect 3185 7642 3191 7644
rect 3247 7642 3271 7644
rect 3327 7642 3351 7644
rect 3407 7642 3431 7644
rect 3487 7642 3493 7644
rect 3247 7590 3249 7642
rect 3429 7590 3431 7642
rect 3185 7588 3191 7590
rect 3247 7588 3271 7590
rect 3327 7588 3351 7590
rect 3407 7588 3431 7590
rect 3487 7588 3493 7590
rect 3185 7579 3493 7588
rect 3792 7472 3844 7478
rect 3792 7414 3844 7420
rect 3516 7404 3568 7410
rect 3516 7346 3568 7352
rect 3332 6928 3384 6934
rect 3332 6870 3384 6876
rect 3344 6798 3372 6870
rect 3528 6798 3556 7346
rect 3608 7268 3660 7274
rect 3608 7210 3660 7216
rect 3620 6866 3648 7210
rect 3700 7200 3752 7206
rect 3700 7142 3752 7148
rect 3608 6860 3660 6866
rect 3608 6802 3660 6808
rect 3332 6792 3384 6798
rect 3332 6734 3384 6740
rect 3516 6792 3568 6798
rect 3516 6734 3568 6740
rect 3056 6724 3108 6730
rect 3056 6666 3108 6672
rect 3516 6656 3568 6662
rect 3516 6598 3568 6604
rect 3185 6556 3493 6565
rect 3185 6554 3191 6556
rect 3247 6554 3271 6556
rect 3327 6554 3351 6556
rect 3407 6554 3431 6556
rect 3487 6554 3493 6556
rect 3247 6502 3249 6554
rect 3429 6502 3431 6554
rect 3185 6500 3191 6502
rect 3247 6500 3271 6502
rect 3327 6500 3351 6502
rect 3407 6500 3431 6502
rect 3487 6500 3493 6502
rect 3185 6491 3493 6500
rect 3056 6384 3108 6390
rect 3056 6326 3108 6332
rect 2964 5772 3016 5778
rect 2964 5714 3016 5720
rect 2872 5704 2924 5710
rect 2872 5646 2924 5652
rect 2884 5302 2912 5646
rect 3068 5370 3096 6326
rect 3424 6248 3476 6254
rect 3424 6190 3476 6196
rect 3436 5778 3464 6190
rect 3528 5914 3556 6598
rect 3620 6118 3648 6802
rect 3712 6186 3740 7142
rect 3804 6798 3832 7414
rect 3976 7404 4028 7410
rect 3976 7346 4028 7352
rect 3884 6928 3936 6934
rect 3988 6882 4016 7346
rect 4448 7002 4476 7754
rect 4436 6996 4488 7002
rect 4436 6938 4488 6944
rect 3936 6876 4016 6882
rect 3884 6870 4016 6876
rect 3896 6854 4016 6870
rect 3988 6798 4016 6854
rect 4068 6860 4120 6866
rect 4068 6802 4120 6808
rect 3792 6792 3844 6798
rect 3792 6734 3844 6740
rect 3976 6792 4028 6798
rect 3976 6734 4028 6740
rect 3884 6656 3936 6662
rect 3884 6598 3936 6604
rect 3896 6322 3924 6598
rect 3884 6316 3936 6322
rect 3884 6258 3936 6264
rect 3988 6202 4016 6734
rect 4080 6458 4108 6802
rect 4344 6724 4396 6730
rect 4344 6666 4396 6672
rect 4160 6656 4212 6662
rect 4160 6598 4212 6604
rect 4068 6452 4120 6458
rect 4068 6394 4120 6400
rect 4172 6322 4200 6598
rect 4356 6458 4384 6666
rect 4344 6452 4396 6458
rect 4344 6394 4396 6400
rect 4160 6316 4212 6322
rect 4160 6258 4212 6264
rect 4252 6248 4304 6254
rect 3988 6196 4252 6202
rect 3988 6190 4304 6196
rect 3700 6180 3752 6186
rect 3988 6174 4292 6190
rect 3700 6122 3752 6128
rect 3608 6112 3660 6118
rect 3608 6054 3660 6060
rect 3516 5908 3568 5914
rect 3516 5850 3568 5856
rect 3424 5772 3476 5778
rect 3424 5714 3476 5720
rect 3712 5710 3740 6122
rect 3976 6112 4028 6118
rect 3976 6054 4028 6060
rect 3988 5710 4016 6054
rect 4080 5846 4108 6174
rect 4448 6066 4476 6938
rect 4540 6390 4568 9302
rect 5368 8974 5396 9318
rect 5676 9276 5984 9285
rect 5676 9274 5682 9276
rect 5738 9274 5762 9276
rect 5818 9274 5842 9276
rect 5898 9274 5922 9276
rect 5978 9274 5984 9276
rect 5738 9222 5740 9274
rect 5920 9222 5922 9274
rect 5676 9220 5682 9222
rect 5738 9220 5762 9222
rect 5818 9220 5842 9222
rect 5898 9220 5922 9222
rect 5978 9220 5984 9222
rect 5676 9211 5984 9220
rect 5448 9104 5500 9110
rect 5448 9046 5500 9052
rect 5460 8974 5488 9046
rect 6564 8974 6592 9551
rect 5356 8968 5408 8974
rect 5356 8910 5408 8916
rect 5448 8968 5500 8974
rect 5448 8910 5500 8916
rect 6552 8968 6604 8974
rect 6552 8910 6604 8916
rect 5172 8900 5224 8906
rect 5172 8842 5224 8848
rect 4712 8288 4764 8294
rect 4712 8230 4764 8236
rect 4724 8090 4752 8230
rect 4712 8084 4764 8090
rect 4712 8026 4764 8032
rect 5184 7886 5212 8842
rect 5368 8498 5396 8910
rect 5356 8492 5408 8498
rect 5356 8434 5408 8440
rect 5460 8378 5488 8910
rect 6336 8732 6644 8741
rect 6336 8730 6342 8732
rect 6398 8730 6422 8732
rect 6478 8730 6502 8732
rect 6558 8730 6582 8732
rect 6638 8730 6644 8732
rect 6398 8678 6400 8730
rect 6580 8678 6582 8730
rect 6336 8676 6342 8678
rect 6398 8676 6422 8678
rect 6478 8676 6502 8678
rect 6558 8676 6582 8678
rect 6638 8676 6644 8678
rect 6336 8667 6644 8676
rect 6748 8634 6776 10610
rect 6828 10600 6880 10606
rect 6828 10542 6880 10548
rect 6840 9042 6868 10542
rect 7116 10062 7144 11698
rect 7104 10056 7156 10062
rect 7104 9998 7156 10004
rect 6828 9036 6880 9042
rect 6828 8978 6880 8984
rect 6920 9036 6972 9042
rect 6920 8978 6972 8984
rect 6736 8628 6788 8634
rect 6736 8570 6788 8576
rect 6748 8514 6776 8570
rect 6656 8486 6776 8514
rect 6840 8498 6868 8978
rect 6828 8492 6880 8498
rect 6656 8430 6684 8486
rect 6828 8434 6880 8440
rect 5368 8350 5488 8378
rect 6644 8424 6696 8430
rect 6644 8366 6696 8372
rect 5368 7886 5396 8350
rect 6736 8288 6788 8294
rect 6736 8230 6788 8236
rect 5676 8188 5984 8197
rect 5676 8186 5682 8188
rect 5738 8186 5762 8188
rect 5818 8186 5842 8188
rect 5898 8186 5922 8188
rect 5978 8186 5984 8188
rect 5738 8134 5740 8186
rect 5920 8134 5922 8186
rect 5676 8132 5682 8134
rect 5738 8132 5762 8134
rect 5818 8132 5842 8134
rect 5898 8132 5922 8134
rect 5978 8132 5984 8134
rect 5676 8123 5984 8132
rect 5172 7880 5224 7886
rect 5172 7822 5224 7828
rect 5356 7880 5408 7886
rect 5356 7822 5408 7828
rect 4712 7744 4764 7750
rect 4712 7686 4764 7692
rect 4620 7200 4672 7206
rect 4620 7142 4672 7148
rect 4528 6384 4580 6390
rect 4528 6326 4580 6332
rect 4632 6322 4660 7142
rect 4724 6458 4752 7686
rect 5184 7546 5212 7822
rect 5908 7744 5960 7750
rect 5908 7686 5960 7692
rect 5172 7540 5224 7546
rect 5172 7482 5224 7488
rect 5920 7478 5948 7686
rect 6336 7644 6644 7653
rect 6336 7642 6342 7644
rect 6398 7642 6422 7644
rect 6478 7642 6502 7644
rect 6558 7642 6582 7644
rect 6638 7642 6644 7644
rect 6398 7590 6400 7642
rect 6580 7590 6582 7642
rect 6336 7588 6342 7590
rect 6398 7588 6422 7590
rect 6478 7588 6502 7590
rect 6558 7588 6582 7590
rect 6638 7588 6644 7590
rect 6336 7579 6644 7588
rect 5908 7472 5960 7478
rect 5908 7414 5960 7420
rect 6644 7472 6696 7478
rect 6644 7414 6696 7420
rect 6184 7336 6236 7342
rect 6184 7278 6236 7284
rect 5676 7100 5984 7109
rect 5676 7098 5682 7100
rect 5738 7098 5762 7100
rect 5818 7098 5842 7100
rect 5898 7098 5922 7100
rect 5978 7098 5984 7100
rect 5738 7046 5740 7098
rect 5920 7046 5922 7098
rect 5676 7044 5682 7046
rect 5738 7044 5762 7046
rect 5818 7044 5842 7046
rect 5898 7044 5922 7046
rect 5978 7044 5984 7046
rect 5676 7035 5984 7044
rect 4896 6860 4948 6866
rect 4896 6802 4948 6808
rect 4712 6452 4764 6458
rect 4712 6394 4764 6400
rect 4620 6316 4672 6322
rect 4620 6258 4672 6264
rect 4264 6038 4476 6066
rect 4068 5840 4120 5846
rect 4068 5782 4120 5788
rect 3700 5704 3752 5710
rect 3700 5646 3752 5652
rect 3976 5704 4028 5710
rect 3976 5646 4028 5652
rect 4264 5642 4292 6038
rect 4908 5914 4936 6802
rect 5816 6656 5868 6662
rect 5816 6598 5868 6604
rect 5828 6322 5856 6598
rect 6092 6384 6144 6390
rect 6092 6326 6144 6332
rect 5816 6316 5868 6322
rect 5816 6258 5868 6264
rect 5676 6012 5984 6021
rect 5676 6010 5682 6012
rect 5738 6010 5762 6012
rect 5818 6010 5842 6012
rect 5898 6010 5922 6012
rect 5978 6010 5984 6012
rect 5738 5958 5740 6010
rect 5920 5958 5922 6010
rect 5676 5956 5682 5958
rect 5738 5956 5762 5958
rect 5818 5956 5842 5958
rect 5898 5956 5922 5958
rect 5978 5956 5984 5958
rect 5676 5947 5984 5956
rect 4896 5908 4948 5914
rect 4896 5850 4948 5856
rect 4252 5636 4304 5642
rect 4252 5578 4304 5584
rect 3185 5468 3493 5477
rect 3185 5466 3191 5468
rect 3247 5466 3271 5468
rect 3327 5466 3351 5468
rect 3407 5466 3431 5468
rect 3487 5466 3493 5468
rect 3247 5414 3249 5466
rect 3429 5414 3431 5466
rect 3185 5412 3191 5414
rect 3247 5412 3271 5414
rect 3327 5412 3351 5414
rect 3407 5412 3431 5414
rect 3487 5412 3493 5414
rect 3185 5403 3493 5412
rect 3056 5364 3108 5370
rect 3056 5306 3108 5312
rect 2872 5296 2924 5302
rect 2872 5238 2924 5244
rect 2136 5228 2188 5234
rect 2136 5170 2188 5176
rect 3608 5228 3660 5234
rect 3608 5170 3660 5176
rect 2525 4924 2833 4933
rect 2525 4922 2531 4924
rect 2587 4922 2611 4924
rect 2667 4922 2691 4924
rect 2747 4922 2771 4924
rect 2827 4922 2833 4924
rect 2587 4870 2589 4922
rect 2769 4870 2771 4922
rect 2525 4868 2531 4870
rect 2587 4868 2611 4870
rect 2667 4868 2691 4870
rect 2747 4868 2771 4870
rect 2827 4868 2833 4870
rect 2525 4859 2833 4868
rect 3620 4758 3648 5170
rect 3976 4820 4028 4826
rect 3976 4762 4028 4768
rect 3608 4752 3660 4758
rect 3608 4694 3660 4700
rect 3185 4380 3493 4389
rect 3185 4378 3191 4380
rect 3247 4378 3271 4380
rect 3327 4378 3351 4380
rect 3407 4378 3431 4380
rect 3487 4378 3493 4380
rect 3247 4326 3249 4378
rect 3429 4326 3431 4378
rect 3185 4324 3191 4326
rect 3247 4324 3271 4326
rect 3327 4324 3351 4326
rect 3407 4324 3431 4326
rect 3487 4324 3493 4326
rect 3185 4315 3493 4324
rect 2525 3836 2833 3845
rect 2525 3834 2531 3836
rect 2587 3834 2611 3836
rect 2667 3834 2691 3836
rect 2747 3834 2771 3836
rect 2827 3834 2833 3836
rect 2587 3782 2589 3834
rect 2769 3782 2771 3834
rect 2525 3780 2531 3782
rect 2587 3780 2611 3782
rect 2667 3780 2691 3782
rect 2747 3780 2771 3782
rect 2827 3780 2833 3782
rect 2525 3771 2833 3780
rect 848 3664 900 3670
rect 846 3632 848 3641
rect 900 3632 902 3641
rect 846 3567 902 3576
rect 3516 3596 3568 3602
rect 3516 3538 3568 3544
rect 3056 3392 3108 3398
rect 3056 3334 3108 3340
rect 3068 2990 3096 3334
rect 3185 3292 3493 3301
rect 3185 3290 3191 3292
rect 3247 3290 3271 3292
rect 3327 3290 3351 3292
rect 3407 3290 3431 3292
rect 3487 3290 3493 3292
rect 3247 3238 3249 3290
rect 3429 3238 3431 3290
rect 3185 3236 3191 3238
rect 3247 3236 3271 3238
rect 3327 3236 3351 3238
rect 3407 3236 3431 3238
rect 3487 3236 3493 3238
rect 3185 3227 3493 3236
rect 3528 3126 3556 3538
rect 3620 3534 3648 4694
rect 3988 3942 4016 4762
rect 4068 4684 4120 4690
rect 4068 4626 4120 4632
rect 3976 3936 4028 3942
rect 3976 3878 4028 3884
rect 4080 3602 4108 4626
rect 4160 4480 4212 4486
rect 4160 4422 4212 4428
rect 4068 3596 4120 3602
rect 4068 3538 4120 3544
rect 3608 3528 3660 3534
rect 3608 3470 3660 3476
rect 3516 3120 3568 3126
rect 3516 3062 3568 3068
rect 848 2984 900 2990
rect 846 2952 848 2961
rect 3056 2984 3108 2990
rect 900 2952 902 2961
rect 3056 2926 3108 2932
rect 846 2887 902 2896
rect 2525 2748 2833 2757
rect 2525 2746 2531 2748
rect 2587 2746 2611 2748
rect 2667 2746 2691 2748
rect 2747 2746 2771 2748
rect 2827 2746 2833 2748
rect 2587 2694 2589 2746
rect 2769 2694 2771 2746
rect 2525 2692 2531 2694
rect 2587 2692 2611 2694
rect 2667 2692 2691 2694
rect 2747 2692 2771 2694
rect 2827 2692 2833 2694
rect 2525 2683 2833 2692
rect 3620 2446 3648 3470
rect 4068 3460 4120 3466
rect 4172 3448 4200 4422
rect 4264 4010 4292 5578
rect 4908 5302 4936 5850
rect 4896 5296 4948 5302
rect 4896 5238 4948 5244
rect 4804 4820 4856 4826
rect 4804 4762 4856 4768
rect 4816 4622 4844 4762
rect 4908 4690 4936 5238
rect 5540 5160 5592 5166
rect 5540 5102 5592 5108
rect 4896 4684 4948 4690
rect 4896 4626 4948 4632
rect 5448 4684 5500 4690
rect 5448 4626 5500 4632
rect 4344 4616 4396 4622
rect 4344 4558 4396 4564
rect 4804 4616 4856 4622
rect 4804 4558 4856 4564
rect 4356 4282 4384 4558
rect 4620 4480 4672 4486
rect 4620 4422 4672 4428
rect 4896 4480 4948 4486
rect 4896 4422 4948 4428
rect 4344 4276 4396 4282
rect 4344 4218 4396 4224
rect 4252 4004 4304 4010
rect 4252 3946 4304 3952
rect 4632 3738 4660 4422
rect 4620 3732 4672 3738
rect 4620 3674 4672 3680
rect 4120 3420 4200 3448
rect 4068 3402 4120 3408
rect 4908 3194 4936 4422
rect 5172 4276 5224 4282
rect 5172 4218 5224 4224
rect 5184 4078 5212 4218
rect 5460 4162 5488 4626
rect 5552 4282 5580 5102
rect 6104 5098 6132 6326
rect 6196 5914 6224 7278
rect 6656 6866 6684 7414
rect 6748 7410 6776 8230
rect 6736 7404 6788 7410
rect 6736 7346 6788 7352
rect 6644 6860 6696 6866
rect 6644 6802 6696 6808
rect 6336 6556 6644 6565
rect 6336 6554 6342 6556
rect 6398 6554 6422 6556
rect 6478 6554 6502 6556
rect 6558 6554 6582 6556
rect 6638 6554 6644 6556
rect 6398 6502 6400 6554
rect 6580 6502 6582 6554
rect 6336 6500 6342 6502
rect 6398 6500 6422 6502
rect 6478 6500 6502 6502
rect 6558 6500 6582 6502
rect 6638 6500 6644 6502
rect 6336 6491 6644 6500
rect 6748 6322 6776 7346
rect 6932 6882 6960 8978
rect 7116 7478 7144 9998
rect 7208 7546 7236 12038
rect 7944 11082 7972 12242
rect 8404 12238 8432 12582
rect 8496 12434 8524 12922
rect 8588 12918 8616 13126
rect 9140 12986 9168 13262
rect 9404 13252 9456 13258
rect 9404 13194 9456 13200
rect 9128 12980 9180 12986
rect 9128 12922 9180 12928
rect 8576 12912 8628 12918
rect 8576 12854 8628 12860
rect 9416 12646 9444 13194
rect 9864 13184 9916 13190
rect 9864 13126 9916 13132
rect 9487 13084 9795 13093
rect 9487 13082 9493 13084
rect 9549 13082 9573 13084
rect 9629 13082 9653 13084
rect 9709 13082 9733 13084
rect 9789 13082 9795 13084
rect 9549 13030 9551 13082
rect 9731 13030 9733 13082
rect 9487 13028 9493 13030
rect 9549 13028 9573 13030
rect 9629 13028 9653 13030
rect 9709 13028 9733 13030
rect 9789 13028 9795 13030
rect 9487 13019 9795 13028
rect 9876 12918 9904 13126
rect 9864 12912 9916 12918
rect 9864 12854 9916 12860
rect 9404 12640 9456 12646
rect 9404 12582 9456 12588
rect 8827 12540 9135 12549
rect 8827 12538 8833 12540
rect 8889 12538 8913 12540
rect 8969 12538 8993 12540
rect 9049 12538 9073 12540
rect 9129 12538 9135 12540
rect 8889 12486 8891 12538
rect 9071 12486 9073 12538
rect 8827 12484 8833 12486
rect 8889 12484 8913 12486
rect 8969 12484 8993 12486
rect 9049 12484 9073 12486
rect 9129 12484 9135 12486
rect 8827 12475 9135 12484
rect 8496 12406 8616 12434
rect 8588 12238 8616 12406
rect 8392 12232 8444 12238
rect 8392 12174 8444 12180
rect 8576 12232 8628 12238
rect 8576 12174 8628 12180
rect 8300 11824 8352 11830
rect 8300 11766 8352 11772
rect 8208 11144 8260 11150
rect 8208 11086 8260 11092
rect 7932 11076 7984 11082
rect 7932 11018 7984 11024
rect 7840 10532 7892 10538
rect 7840 10474 7892 10480
rect 7656 8628 7708 8634
rect 7656 8570 7708 8576
rect 7668 8537 7696 8570
rect 7654 8528 7710 8537
rect 7654 8463 7710 8472
rect 7288 8288 7340 8294
rect 7288 8230 7340 8236
rect 7300 7750 7328 8230
rect 7668 7886 7696 8463
rect 7852 8430 7880 10474
rect 7944 9586 7972 11018
rect 8116 10668 8168 10674
rect 8116 10610 8168 10616
rect 8128 10470 8156 10610
rect 8220 10470 8248 11086
rect 8116 10464 8168 10470
rect 8116 10406 8168 10412
rect 8208 10464 8260 10470
rect 8208 10406 8260 10412
rect 8128 10044 8156 10406
rect 8208 10056 8260 10062
rect 8128 10016 8208 10044
rect 8208 9998 8260 10004
rect 8116 9920 8168 9926
rect 8116 9862 8168 9868
rect 8128 9654 8156 9862
rect 8312 9738 8340 11766
rect 8404 11098 8432 12174
rect 8404 11070 8524 11098
rect 8392 11008 8444 11014
rect 8392 10950 8444 10956
rect 8404 10810 8432 10950
rect 8392 10804 8444 10810
rect 8392 10746 8444 10752
rect 8404 10198 8432 10746
rect 8496 10538 8524 11070
rect 8588 10674 8616 12174
rect 9416 12102 9444 12582
rect 10244 12306 10272 13806
rect 13372 13705 13400 13806
rect 13358 13696 13414 13705
rect 11978 13628 12286 13637
rect 13358 13631 13414 13640
rect 11978 13626 11984 13628
rect 12040 13626 12064 13628
rect 12120 13626 12144 13628
rect 12200 13626 12224 13628
rect 12280 13626 12286 13628
rect 12040 13574 12042 13626
rect 12222 13574 12224 13626
rect 11978 13572 11984 13574
rect 12040 13572 12064 13574
rect 12120 13572 12144 13574
rect 12200 13572 12224 13574
rect 12280 13572 12286 13574
rect 11978 13563 12286 13572
rect 10416 13320 10468 13326
rect 10416 13262 10468 13268
rect 10428 12850 10456 13262
rect 13360 13184 13412 13190
rect 13360 13126 13412 13132
rect 12638 13084 12946 13093
rect 12638 13082 12644 13084
rect 12700 13082 12724 13084
rect 12780 13082 12804 13084
rect 12860 13082 12884 13084
rect 12940 13082 12946 13084
rect 12700 13030 12702 13082
rect 12882 13030 12884 13082
rect 12638 13028 12644 13030
rect 12700 13028 12724 13030
rect 12780 13028 12804 13030
rect 12860 13028 12884 13030
rect 12940 13028 12946 13030
rect 12638 13019 12946 13028
rect 13372 13025 13400 13126
rect 13358 13016 13414 13025
rect 13358 12951 13414 12960
rect 10416 12844 10468 12850
rect 10416 12786 10468 12792
rect 10324 12640 10376 12646
rect 10324 12582 10376 12588
rect 10232 12300 10284 12306
rect 10232 12242 10284 12248
rect 9864 12164 9916 12170
rect 9864 12106 9916 12112
rect 9404 12096 9456 12102
rect 9404 12038 9456 12044
rect 8827 11452 9135 11461
rect 8827 11450 8833 11452
rect 8889 11450 8913 11452
rect 8969 11450 8993 11452
rect 9049 11450 9073 11452
rect 9129 11450 9135 11452
rect 8889 11398 8891 11450
rect 9071 11398 9073 11450
rect 8827 11396 8833 11398
rect 8889 11396 8913 11398
rect 8969 11396 8993 11398
rect 9049 11396 9073 11398
rect 9129 11396 9135 11398
rect 8827 11387 9135 11396
rect 9416 11354 9444 12038
rect 9487 11996 9795 12005
rect 9487 11994 9493 11996
rect 9549 11994 9573 11996
rect 9629 11994 9653 11996
rect 9709 11994 9733 11996
rect 9789 11994 9795 11996
rect 9549 11942 9551 11994
rect 9731 11942 9733 11994
rect 9487 11940 9493 11942
rect 9549 11940 9573 11942
rect 9629 11940 9653 11942
rect 9709 11940 9733 11942
rect 9789 11940 9795 11942
rect 9487 11931 9795 11940
rect 9876 11354 9904 12106
rect 10244 11898 10272 12242
rect 10336 12170 10364 12582
rect 10324 12164 10376 12170
rect 10324 12106 10376 12112
rect 10232 11892 10284 11898
rect 10232 11834 10284 11840
rect 9404 11348 9456 11354
rect 9404 11290 9456 11296
rect 9864 11348 9916 11354
rect 9864 11290 9916 11296
rect 9220 11076 9272 11082
rect 9220 11018 9272 11024
rect 8576 10668 8628 10674
rect 8576 10610 8628 10616
rect 9232 10538 9260 11018
rect 9416 10810 9444 11290
rect 9956 11008 10008 11014
rect 9956 10950 10008 10956
rect 9487 10908 9795 10917
rect 9487 10906 9493 10908
rect 9549 10906 9573 10908
rect 9629 10906 9653 10908
rect 9709 10906 9733 10908
rect 9789 10906 9795 10908
rect 9549 10854 9551 10906
rect 9731 10854 9733 10906
rect 9487 10852 9493 10854
rect 9549 10852 9573 10854
rect 9629 10852 9653 10854
rect 9709 10852 9733 10854
rect 9789 10852 9795 10854
rect 9487 10843 9795 10852
rect 9404 10804 9456 10810
rect 9404 10746 9456 10752
rect 9588 10804 9640 10810
rect 9588 10746 9640 10752
rect 9324 10674 9536 10690
rect 9312 10668 9536 10674
rect 9364 10662 9536 10668
rect 9312 10610 9364 10616
rect 9508 10606 9536 10662
rect 9600 10606 9628 10746
rect 9680 10736 9732 10742
rect 9680 10678 9732 10684
rect 9496 10600 9548 10606
rect 9496 10542 9548 10548
rect 9588 10600 9640 10606
rect 9588 10542 9640 10548
rect 8484 10532 8536 10538
rect 8484 10474 8536 10480
rect 9220 10532 9272 10538
rect 9220 10474 9272 10480
rect 8576 10464 8628 10470
rect 8576 10406 8628 10412
rect 9232 10418 9260 10474
rect 8392 10192 8444 10198
rect 8392 10134 8444 10140
rect 8484 10056 8536 10062
rect 8484 9998 8536 10004
rect 8392 9920 8444 9926
rect 8392 9862 8444 9868
rect 8220 9710 8340 9738
rect 8116 9648 8168 9654
rect 8116 9590 8168 9596
rect 7932 9580 7984 9586
rect 7932 9522 7984 9528
rect 8220 9042 8248 9710
rect 8404 9178 8432 9862
rect 8496 9722 8524 9998
rect 8484 9716 8536 9722
rect 8484 9658 8536 9664
rect 8392 9172 8444 9178
rect 8392 9114 8444 9120
rect 8208 9036 8260 9042
rect 8208 8978 8260 8984
rect 8392 8832 8444 8838
rect 8392 8774 8444 8780
rect 8300 8628 8352 8634
rect 8300 8570 8352 8576
rect 7932 8560 7984 8566
rect 8312 8514 8340 8570
rect 7984 8508 8340 8514
rect 7932 8502 8340 8508
rect 7944 8486 8340 8502
rect 8404 8498 8432 8774
rect 8496 8634 8524 9658
rect 8588 9178 8616 10406
rect 9232 10390 9352 10418
rect 8827 10364 9135 10373
rect 8827 10362 8833 10364
rect 8889 10362 8913 10364
rect 8969 10362 8993 10364
rect 9049 10362 9073 10364
rect 9129 10362 9135 10364
rect 8889 10310 8891 10362
rect 9071 10310 9073 10362
rect 8827 10308 8833 10310
rect 8889 10308 8913 10310
rect 8969 10308 8993 10310
rect 9049 10308 9073 10310
rect 9129 10308 9135 10310
rect 8827 10299 9135 10308
rect 9220 9988 9272 9994
rect 9220 9930 9272 9936
rect 8668 9920 8720 9926
rect 8668 9862 8720 9868
rect 8576 9172 8628 9178
rect 8576 9114 8628 9120
rect 8576 8968 8628 8974
rect 8576 8910 8628 8916
rect 8484 8628 8536 8634
rect 8484 8570 8536 8576
rect 8392 8492 8444 8498
rect 8392 8434 8444 8440
rect 7840 8424 7892 8430
rect 7840 8366 7892 8372
rect 8484 8424 8536 8430
rect 8484 8366 8536 8372
rect 8392 8356 8444 8362
rect 8392 8298 8444 8304
rect 7656 7880 7708 7886
rect 7656 7822 7708 7828
rect 8300 7880 8352 7886
rect 8300 7822 8352 7828
rect 7288 7744 7340 7750
rect 7288 7686 7340 7692
rect 7196 7540 7248 7546
rect 7196 7482 7248 7488
rect 7104 7472 7156 7478
rect 7104 7414 7156 7420
rect 7380 7404 7432 7410
rect 7380 7346 7432 7352
rect 6840 6854 6960 6882
rect 6736 6316 6788 6322
rect 6736 6258 6788 6264
rect 6184 5908 6236 5914
rect 6184 5850 6236 5856
rect 6336 5468 6644 5477
rect 6336 5466 6342 5468
rect 6398 5466 6422 5468
rect 6478 5466 6502 5468
rect 6558 5466 6582 5468
rect 6638 5466 6644 5468
rect 6398 5414 6400 5466
rect 6580 5414 6582 5466
rect 6336 5412 6342 5414
rect 6398 5412 6422 5414
rect 6478 5412 6502 5414
rect 6558 5412 6582 5414
rect 6638 5412 6644 5414
rect 6336 5403 6644 5412
rect 6092 5092 6144 5098
rect 6092 5034 6144 5040
rect 6000 5024 6052 5030
rect 6000 4966 6052 4972
rect 5676 4924 5984 4933
rect 5676 4922 5682 4924
rect 5738 4922 5762 4924
rect 5818 4922 5842 4924
rect 5898 4922 5922 4924
rect 5978 4922 5984 4924
rect 5738 4870 5740 4922
rect 5920 4870 5922 4922
rect 5676 4868 5682 4870
rect 5738 4868 5762 4870
rect 5818 4868 5842 4870
rect 5898 4868 5922 4870
rect 5978 4868 5984 4870
rect 5676 4859 5984 4868
rect 5632 4548 5684 4554
rect 5632 4490 5684 4496
rect 5724 4548 5776 4554
rect 5724 4490 5776 4496
rect 5540 4276 5592 4282
rect 5540 4218 5592 4224
rect 5264 4140 5316 4146
rect 5460 4134 5580 4162
rect 5264 4082 5316 4088
rect 5172 4072 5224 4078
rect 5172 4014 5224 4020
rect 4988 4004 5040 4010
rect 4988 3946 5040 3952
rect 4896 3188 4948 3194
rect 4896 3130 4948 3136
rect 4160 3120 4212 3126
rect 4160 3062 4212 3068
rect 4172 2650 4200 3062
rect 5000 2990 5028 3946
rect 5184 3194 5212 4014
rect 5276 3738 5304 4082
rect 5448 4072 5500 4078
rect 5448 4014 5500 4020
rect 5264 3732 5316 3738
rect 5264 3674 5316 3680
rect 5172 3188 5224 3194
rect 5172 3130 5224 3136
rect 5460 3058 5488 4014
rect 5552 3602 5580 4134
rect 5644 4010 5672 4490
rect 5736 4282 5764 4490
rect 5724 4276 5776 4282
rect 5724 4218 5776 4224
rect 6012 4146 6040 4966
rect 6092 4480 6144 4486
rect 6092 4422 6144 4428
rect 6000 4140 6052 4146
rect 6000 4082 6052 4088
rect 5632 4004 5684 4010
rect 5632 3946 5684 3952
rect 6000 3936 6052 3942
rect 6000 3878 6052 3884
rect 5676 3836 5984 3845
rect 5676 3834 5682 3836
rect 5738 3834 5762 3836
rect 5818 3834 5842 3836
rect 5898 3834 5922 3836
rect 5978 3834 5984 3836
rect 5738 3782 5740 3834
rect 5920 3782 5922 3834
rect 5676 3780 5682 3782
rect 5738 3780 5762 3782
rect 5818 3780 5842 3782
rect 5898 3780 5922 3782
rect 5978 3780 5984 3782
rect 5676 3771 5984 3780
rect 6012 3618 6040 3878
rect 5540 3596 5592 3602
rect 5540 3538 5592 3544
rect 5828 3590 6040 3618
rect 5828 3534 5856 3590
rect 5816 3528 5868 3534
rect 5816 3470 5868 3476
rect 6104 3194 6132 4422
rect 6336 4380 6644 4389
rect 6336 4378 6342 4380
rect 6398 4378 6422 4380
rect 6478 4378 6502 4380
rect 6558 4378 6582 4380
rect 6638 4378 6644 4380
rect 6398 4326 6400 4378
rect 6580 4326 6582 4378
rect 6336 4324 6342 4326
rect 6398 4324 6422 4326
rect 6478 4324 6502 4326
rect 6558 4324 6582 4326
rect 6638 4324 6644 4326
rect 6336 4315 6644 4324
rect 6184 4208 6236 4214
rect 6184 4150 6236 4156
rect 6196 3194 6224 4150
rect 6748 4010 6776 6258
rect 6840 5710 6868 6854
rect 7392 6730 7420 7346
rect 8312 6934 8340 7822
rect 8300 6928 8352 6934
rect 8300 6870 8352 6876
rect 7380 6724 7432 6730
rect 7380 6666 7432 6672
rect 8300 6724 8352 6730
rect 8300 6666 8352 6672
rect 7392 6322 7420 6666
rect 8312 6458 8340 6666
rect 8300 6452 8352 6458
rect 8300 6394 8352 6400
rect 7380 6316 7432 6322
rect 7380 6258 7432 6264
rect 6828 5704 6880 5710
rect 6828 5646 6880 5652
rect 6828 4752 6880 4758
rect 6828 4694 6880 4700
rect 6840 4146 6868 4694
rect 6828 4140 6880 4146
rect 6828 4082 6880 4088
rect 6736 4004 6788 4010
rect 6736 3946 6788 3952
rect 6336 3292 6644 3301
rect 6336 3290 6342 3292
rect 6398 3290 6422 3292
rect 6478 3290 6502 3292
rect 6558 3290 6582 3292
rect 6638 3290 6644 3292
rect 6398 3238 6400 3290
rect 6580 3238 6582 3290
rect 6336 3236 6342 3238
rect 6398 3236 6422 3238
rect 6478 3236 6502 3238
rect 6558 3236 6582 3238
rect 6638 3236 6644 3238
rect 6336 3227 6644 3236
rect 6092 3188 6144 3194
rect 6092 3130 6144 3136
rect 6184 3188 6236 3194
rect 6184 3130 6236 3136
rect 6840 3058 6868 4082
rect 6920 3460 6972 3466
rect 6920 3402 6972 3408
rect 6932 3194 6960 3402
rect 6920 3188 6972 3194
rect 6920 3130 6972 3136
rect 5448 3052 5500 3058
rect 5448 2994 5500 3000
rect 6828 3052 6880 3058
rect 6828 2994 6880 3000
rect 4988 2984 5040 2990
rect 4988 2926 5040 2932
rect 5676 2748 5984 2757
rect 5676 2746 5682 2748
rect 5738 2746 5762 2748
rect 5818 2746 5842 2748
rect 5898 2746 5922 2748
rect 5978 2746 5984 2748
rect 5738 2694 5740 2746
rect 5920 2694 5922 2746
rect 5676 2692 5682 2694
rect 5738 2692 5762 2694
rect 5818 2692 5842 2694
rect 5898 2692 5922 2694
rect 5978 2692 5984 2694
rect 5676 2683 5984 2692
rect 7392 2650 7420 6258
rect 8404 6254 8432 8298
rect 8496 8022 8524 8366
rect 8484 8016 8536 8022
rect 8484 7958 8536 7964
rect 8484 7744 8536 7750
rect 8484 7686 8536 7692
rect 7932 6248 7984 6254
rect 7932 6190 7984 6196
rect 8392 6248 8444 6254
rect 8392 6190 8444 6196
rect 8496 6202 8524 7686
rect 8588 7546 8616 8910
rect 8680 8634 8708 9862
rect 9128 9716 9180 9722
rect 9128 9658 9180 9664
rect 9140 9364 9168 9658
rect 9232 9654 9260 9930
rect 9324 9926 9352 10390
rect 9404 10260 9456 10266
rect 9404 10202 9456 10208
rect 9312 9920 9364 9926
rect 9312 9862 9364 9868
rect 9220 9648 9272 9654
rect 9220 9590 9272 9596
rect 9140 9336 9260 9364
rect 8827 9276 9135 9285
rect 8827 9274 8833 9276
rect 8889 9274 8913 9276
rect 8969 9274 8993 9276
rect 9049 9274 9073 9276
rect 9129 9274 9135 9276
rect 8889 9222 8891 9274
rect 9071 9222 9073 9274
rect 8827 9220 8833 9222
rect 8889 9220 8913 9222
rect 8969 9220 8993 9222
rect 9049 9220 9073 9222
rect 9129 9220 9135 9222
rect 8827 9211 9135 9220
rect 8668 8628 8720 8634
rect 8668 8570 8720 8576
rect 9232 8566 9260 9336
rect 9416 8906 9444 10202
rect 9692 10198 9720 10678
rect 9968 10674 9996 10950
rect 9956 10668 10008 10674
rect 9956 10610 10008 10616
rect 10324 10668 10376 10674
rect 10324 10610 10376 10616
rect 9680 10192 9732 10198
rect 9680 10134 9732 10140
rect 9968 10130 9996 10610
rect 9956 10124 10008 10130
rect 9956 10066 10008 10072
rect 9487 9820 9795 9829
rect 9487 9818 9493 9820
rect 9549 9818 9573 9820
rect 9629 9818 9653 9820
rect 9709 9818 9733 9820
rect 9789 9818 9795 9820
rect 9549 9766 9551 9818
rect 9731 9766 9733 9818
rect 9487 9764 9493 9766
rect 9549 9764 9573 9766
rect 9629 9764 9653 9766
rect 9709 9764 9733 9766
rect 9789 9764 9795 9766
rect 9487 9755 9795 9764
rect 9968 9722 9996 10066
rect 9956 9716 10008 9722
rect 9956 9658 10008 9664
rect 10336 8974 10364 10610
rect 10428 9926 10456 12786
rect 12440 12640 12492 12646
rect 12440 12582 12492 12588
rect 11978 12540 12286 12549
rect 11978 12538 11984 12540
rect 12040 12538 12064 12540
rect 12120 12538 12144 12540
rect 12200 12538 12224 12540
rect 12280 12538 12286 12540
rect 12040 12486 12042 12538
rect 12222 12486 12224 12538
rect 11978 12484 11984 12486
rect 12040 12484 12064 12486
rect 12120 12484 12144 12486
rect 12200 12484 12224 12486
rect 12280 12484 12286 12486
rect 11978 12475 12286 12484
rect 11520 12300 11572 12306
rect 11520 12242 11572 12248
rect 11428 12164 11480 12170
rect 11428 12106 11480 12112
rect 10876 12096 10928 12102
rect 10876 12038 10928 12044
rect 10784 11892 10836 11898
rect 10784 11834 10836 11840
rect 10600 11688 10652 11694
rect 10600 11630 10652 11636
rect 10612 11150 10640 11630
rect 10796 11150 10824 11834
rect 10888 11150 10916 12038
rect 11440 11898 11468 12106
rect 11428 11892 11480 11898
rect 11428 11834 11480 11840
rect 10968 11824 11020 11830
rect 10968 11766 11020 11772
rect 10980 11286 11008 11766
rect 11060 11756 11112 11762
rect 11060 11698 11112 11704
rect 10968 11280 11020 11286
rect 10968 11222 11020 11228
rect 10508 11144 10560 11150
rect 10508 11086 10560 11092
rect 10600 11144 10652 11150
rect 10600 11086 10652 11092
rect 10784 11144 10836 11150
rect 10784 11086 10836 11092
rect 10876 11144 10928 11150
rect 10876 11086 10928 11092
rect 10416 9920 10468 9926
rect 10416 9862 10468 9868
rect 10520 9722 10548 11086
rect 10612 10742 10640 11086
rect 10600 10736 10652 10742
rect 10600 10678 10652 10684
rect 10796 10674 10824 11086
rect 10888 10810 10916 11086
rect 11072 11082 11100 11698
rect 11428 11212 11480 11218
rect 11428 11154 11480 11160
rect 11060 11076 11112 11082
rect 11060 11018 11112 11024
rect 11152 11008 11204 11014
rect 11152 10950 11204 10956
rect 10876 10804 10928 10810
rect 10876 10746 10928 10752
rect 11164 10674 11192 10950
rect 11440 10810 11468 11154
rect 11428 10804 11480 10810
rect 11428 10746 11480 10752
rect 11532 10674 11560 12242
rect 12452 12170 12480 12582
rect 12440 12164 12492 12170
rect 12440 12106 12492 12112
rect 12992 12096 13044 12102
rect 12992 12038 13044 12044
rect 12638 11996 12946 12005
rect 12638 11994 12644 11996
rect 12700 11994 12724 11996
rect 12780 11994 12804 11996
rect 12860 11994 12884 11996
rect 12940 11994 12946 11996
rect 12700 11942 12702 11994
rect 12882 11942 12884 11994
rect 12638 11940 12644 11942
rect 12700 11940 12724 11942
rect 12780 11940 12804 11942
rect 12860 11940 12884 11942
rect 12940 11940 12946 11942
rect 12638 11931 12946 11940
rect 11704 11756 11756 11762
rect 11704 11698 11756 11704
rect 12348 11756 12400 11762
rect 12348 11698 12400 11704
rect 11716 11354 11744 11698
rect 11978 11452 12286 11461
rect 11978 11450 11984 11452
rect 12040 11450 12064 11452
rect 12120 11450 12144 11452
rect 12200 11450 12224 11452
rect 12280 11450 12286 11452
rect 12040 11398 12042 11450
rect 12222 11398 12224 11450
rect 11978 11396 11984 11398
rect 12040 11396 12064 11398
rect 12120 11396 12144 11398
rect 12200 11396 12224 11398
rect 12280 11396 12286 11398
rect 11978 11387 12286 11396
rect 12360 11354 12388 11698
rect 11704 11348 11756 11354
rect 11704 11290 11756 11296
rect 12348 11348 12400 11354
rect 12348 11290 12400 11296
rect 12256 11280 12308 11286
rect 12256 11222 12308 11228
rect 11612 11212 11664 11218
rect 11612 11154 11664 11160
rect 12072 11212 12124 11218
rect 12072 11154 12124 11160
rect 10784 10668 10836 10674
rect 10784 10610 10836 10616
rect 11152 10668 11204 10674
rect 11152 10610 11204 10616
rect 11520 10668 11572 10674
rect 11520 10610 11572 10616
rect 11244 10600 11296 10606
rect 11244 10542 11296 10548
rect 11060 10464 11112 10470
rect 11060 10406 11112 10412
rect 11072 9926 11100 10406
rect 11256 10266 11284 10542
rect 11244 10260 11296 10266
rect 11244 10202 11296 10208
rect 11428 10056 11480 10062
rect 11428 9998 11480 10004
rect 11440 9926 11468 9998
rect 11060 9920 11112 9926
rect 11060 9862 11112 9868
rect 11336 9920 11388 9926
rect 11336 9862 11388 9868
rect 11428 9920 11480 9926
rect 11428 9862 11480 9868
rect 10508 9716 10560 9722
rect 10508 9658 10560 9664
rect 11072 9674 11100 9862
rect 11072 9646 11192 9674
rect 11060 9512 11112 9518
rect 11060 9454 11112 9460
rect 11072 9178 11100 9454
rect 11060 9172 11112 9178
rect 11060 9114 11112 9120
rect 11164 9058 11192 9646
rect 11348 9110 11376 9862
rect 11532 9586 11560 10610
rect 11624 9722 11652 11154
rect 11796 11144 11848 11150
rect 12084 11098 12112 11154
rect 12268 11150 12296 11222
rect 13004 11218 13032 12038
rect 12992 11212 13044 11218
rect 12992 11154 13044 11160
rect 11796 11086 11848 11092
rect 11704 10804 11756 10810
rect 11704 10746 11756 10752
rect 11716 10062 11744 10746
rect 11808 10198 11836 11086
rect 11900 11082 12112 11098
rect 12256 11144 12308 11150
rect 12256 11086 12308 11092
rect 11900 11076 12124 11082
rect 11900 11070 12072 11076
rect 11796 10192 11848 10198
rect 11796 10134 11848 10140
rect 11704 10056 11756 10062
rect 11704 9998 11756 10004
rect 11612 9716 11664 9722
rect 11612 9658 11664 9664
rect 11520 9580 11572 9586
rect 11520 9522 11572 9528
rect 11072 9030 11192 9058
rect 11336 9104 11388 9110
rect 11336 9046 11388 9052
rect 11624 9042 11652 9658
rect 11612 9036 11664 9042
rect 10324 8968 10376 8974
rect 10324 8910 10376 8916
rect 10784 8968 10836 8974
rect 10784 8910 10836 8916
rect 9404 8900 9456 8906
rect 9404 8842 9456 8848
rect 10048 8900 10100 8906
rect 10048 8842 10100 8848
rect 9487 8732 9795 8741
rect 9487 8730 9493 8732
rect 9549 8730 9573 8732
rect 9629 8730 9653 8732
rect 9709 8730 9733 8732
rect 9789 8730 9795 8732
rect 9549 8678 9551 8730
rect 9731 8678 9733 8730
rect 9487 8676 9493 8678
rect 9549 8676 9573 8678
rect 9629 8676 9653 8678
rect 9709 8676 9733 8678
rect 9789 8676 9795 8678
rect 9487 8667 9795 8676
rect 9220 8560 9272 8566
rect 8666 8528 8722 8537
rect 9220 8502 9272 8508
rect 8666 8463 8668 8472
rect 8720 8463 8722 8472
rect 8668 8434 8720 8440
rect 8668 8288 8720 8294
rect 8668 8230 8720 8236
rect 8576 7540 8628 7546
rect 8576 7482 8628 7488
rect 8576 7404 8628 7410
rect 8576 7346 8628 7352
rect 8588 6361 8616 7346
rect 8680 7342 8708 8230
rect 8827 8188 9135 8197
rect 8827 8186 8833 8188
rect 8889 8186 8913 8188
rect 8969 8186 8993 8188
rect 9049 8186 9073 8188
rect 9129 8186 9135 8188
rect 8889 8134 8891 8186
rect 9071 8134 9073 8186
rect 8827 8132 8833 8134
rect 8889 8132 8913 8134
rect 8969 8132 8993 8134
rect 9049 8132 9073 8134
rect 9129 8132 9135 8134
rect 8827 8123 9135 8132
rect 10060 7886 10088 8842
rect 10140 8288 10192 8294
rect 10140 8230 10192 8236
rect 10152 8022 10180 8230
rect 10140 8016 10192 8022
rect 10140 7958 10192 7964
rect 8760 7880 8812 7886
rect 8760 7822 8812 7828
rect 9956 7880 10008 7886
rect 9956 7822 10008 7828
rect 10048 7880 10100 7886
rect 10048 7822 10100 7828
rect 8668 7336 8720 7342
rect 8668 7278 8720 7284
rect 8772 7188 8800 7822
rect 9864 7744 9916 7750
rect 9864 7686 9916 7692
rect 9487 7644 9795 7653
rect 9487 7642 9493 7644
rect 9549 7642 9573 7644
rect 9629 7642 9653 7644
rect 9709 7642 9733 7644
rect 9789 7642 9795 7644
rect 9549 7590 9551 7642
rect 9731 7590 9733 7642
rect 9487 7588 9493 7590
rect 9549 7588 9573 7590
rect 9629 7588 9653 7590
rect 9709 7588 9733 7590
rect 9789 7588 9795 7590
rect 9487 7579 9795 7588
rect 8852 7540 8904 7546
rect 8852 7482 8904 7488
rect 8864 7206 8892 7482
rect 9876 7478 9904 7686
rect 9968 7562 9996 7822
rect 9968 7546 10088 7562
rect 9956 7540 10088 7546
rect 10008 7534 10088 7540
rect 9956 7482 10008 7488
rect 9864 7472 9916 7478
rect 9864 7414 9916 7420
rect 9404 7404 9456 7410
rect 9404 7346 9456 7352
rect 8680 7160 8800 7188
rect 8852 7200 8904 7206
rect 8574 6352 8630 6361
rect 8574 6287 8630 6296
rect 7944 4826 7972 6190
rect 8496 6174 8616 6202
rect 8680 6186 8708 7160
rect 8852 7142 8904 7148
rect 8827 7100 9135 7109
rect 8827 7098 8833 7100
rect 8889 7098 8913 7100
rect 8969 7098 8993 7100
rect 9049 7098 9073 7100
rect 9129 7098 9135 7100
rect 8889 7046 8891 7098
rect 9071 7046 9073 7098
rect 8827 7044 8833 7046
rect 8889 7044 8913 7046
rect 8969 7044 8993 7046
rect 9049 7044 9073 7046
rect 9129 7044 9135 7046
rect 8827 7035 9135 7044
rect 9312 6996 9364 7002
rect 9312 6938 9364 6944
rect 8852 6928 8904 6934
rect 8852 6870 8904 6876
rect 9220 6928 9272 6934
rect 9220 6870 9272 6876
rect 8864 6322 8892 6870
rect 9232 6798 9260 6870
rect 9220 6792 9272 6798
rect 9220 6734 9272 6740
rect 9036 6656 9088 6662
rect 9036 6598 9088 6604
rect 9048 6458 9076 6598
rect 9324 6458 9352 6938
rect 9036 6452 9088 6458
rect 9036 6394 9088 6400
rect 9312 6452 9364 6458
rect 9312 6394 9364 6400
rect 9416 6390 9444 7346
rect 9496 7336 9548 7342
rect 9496 7278 9548 7284
rect 9508 6866 9536 7278
rect 9680 6996 9732 7002
rect 9680 6938 9732 6944
rect 9496 6860 9548 6866
rect 9496 6802 9548 6808
rect 9692 6662 9720 6938
rect 10060 6798 10088 7534
rect 10152 6798 10180 7958
rect 10336 7886 10364 8910
rect 10600 8560 10652 8566
rect 10600 8502 10652 8508
rect 10612 7954 10640 8502
rect 10796 8294 10824 8910
rect 10876 8492 10928 8498
rect 10876 8434 10928 8440
rect 10784 8288 10836 8294
rect 10784 8230 10836 8236
rect 10600 7948 10652 7954
rect 10600 7890 10652 7896
rect 10888 7886 10916 8434
rect 11072 7886 11100 9030
rect 11612 8978 11664 8984
rect 11336 8560 11388 8566
rect 11336 8502 11388 8508
rect 11152 7948 11204 7954
rect 11152 7890 11204 7896
rect 10324 7880 10376 7886
rect 10324 7822 10376 7828
rect 10876 7880 10928 7886
rect 10876 7822 10928 7828
rect 11060 7880 11112 7886
rect 11060 7822 11112 7828
rect 10336 7002 10364 7822
rect 10784 7744 10836 7750
rect 10784 7686 10836 7692
rect 10796 7342 10824 7686
rect 10888 7562 10916 7822
rect 11072 7750 11100 7822
rect 11060 7744 11112 7750
rect 11060 7686 11112 7692
rect 10888 7546 11100 7562
rect 10888 7540 11112 7546
rect 10888 7534 11060 7540
rect 10784 7336 10836 7342
rect 10784 7278 10836 7284
rect 10508 7200 10560 7206
rect 10508 7142 10560 7148
rect 10324 6996 10376 7002
rect 10324 6938 10376 6944
rect 10416 6860 10468 6866
rect 10416 6802 10468 6808
rect 10048 6792 10100 6798
rect 10048 6734 10100 6740
rect 10140 6792 10192 6798
rect 10140 6734 10192 6740
rect 10232 6792 10284 6798
rect 10232 6734 10284 6740
rect 9680 6656 9732 6662
rect 9680 6598 9732 6604
rect 9864 6656 9916 6662
rect 9864 6598 9916 6604
rect 10048 6656 10100 6662
rect 10048 6598 10100 6604
rect 9487 6556 9795 6565
rect 9487 6554 9493 6556
rect 9549 6554 9573 6556
rect 9629 6554 9653 6556
rect 9709 6554 9733 6556
rect 9789 6554 9795 6556
rect 9549 6502 9551 6554
rect 9731 6502 9733 6554
rect 9487 6500 9493 6502
rect 9549 6500 9573 6502
rect 9629 6500 9653 6502
rect 9709 6500 9733 6502
rect 9789 6500 9795 6502
rect 9487 6491 9795 6500
rect 9876 6458 9904 6598
rect 9864 6452 9916 6458
rect 9692 6412 9864 6440
rect 9404 6384 9456 6390
rect 9404 6326 9456 6332
rect 9586 6352 9642 6361
rect 8852 6316 8904 6322
rect 9692 6322 9720 6412
rect 9864 6394 9916 6400
rect 10060 6322 10088 6598
rect 10244 6390 10272 6734
rect 10232 6384 10284 6390
rect 10232 6326 10284 6332
rect 9586 6287 9588 6296
rect 8852 6258 8904 6264
rect 9640 6287 9642 6296
rect 9680 6316 9732 6322
rect 9588 6258 9640 6264
rect 9680 6258 9732 6264
rect 10048 6316 10100 6322
rect 10048 6258 10100 6264
rect 8864 6225 8892 6258
rect 9312 6248 9364 6254
rect 8850 6216 8906 6225
rect 8484 6112 8536 6118
rect 8484 6054 8536 6060
rect 7932 4820 7984 4826
rect 7932 4762 7984 4768
rect 7656 4072 7708 4078
rect 7656 4014 7708 4020
rect 7668 3738 7696 4014
rect 7656 3732 7708 3738
rect 7656 3674 7708 3680
rect 7944 3534 7972 4762
rect 8300 4548 8352 4554
rect 8300 4490 8352 4496
rect 8312 3942 8340 4490
rect 8392 4140 8444 4146
rect 8392 4082 8444 4088
rect 8300 3936 8352 3942
rect 8300 3878 8352 3884
rect 7932 3528 7984 3534
rect 7932 3470 7984 3476
rect 7944 3058 7972 3470
rect 8404 3194 8432 4082
rect 8496 3602 8524 6054
rect 8588 4690 8616 6174
rect 8668 6180 8720 6186
rect 9312 6190 9364 6196
rect 8850 6151 8906 6160
rect 8668 6122 8720 6128
rect 8827 6012 9135 6021
rect 8827 6010 8833 6012
rect 8889 6010 8913 6012
rect 8969 6010 8993 6012
rect 9049 6010 9073 6012
rect 9129 6010 9135 6012
rect 8889 5958 8891 6010
rect 9071 5958 9073 6010
rect 8827 5956 8833 5958
rect 8889 5956 8913 5958
rect 8969 5956 8993 5958
rect 9049 5956 9073 5958
rect 9129 5956 9135 5958
rect 8827 5947 9135 5956
rect 8827 4924 9135 4933
rect 8827 4922 8833 4924
rect 8889 4922 8913 4924
rect 8969 4922 8993 4924
rect 9049 4922 9073 4924
rect 9129 4922 9135 4924
rect 8889 4870 8891 4922
rect 9071 4870 9073 4922
rect 8827 4868 8833 4870
rect 8889 4868 8913 4870
rect 8969 4868 8993 4870
rect 9049 4868 9073 4870
rect 9129 4868 9135 4870
rect 8827 4859 9135 4868
rect 8576 4684 8628 4690
rect 8576 4626 8628 4632
rect 9324 4622 9352 6190
rect 9600 6118 9628 6258
rect 10244 6225 10272 6326
rect 10230 6216 10286 6225
rect 10230 6151 10286 6160
rect 10428 6202 10456 6802
rect 10520 6390 10548 7142
rect 10692 6928 10744 6934
rect 10692 6870 10744 6876
rect 10600 6656 10652 6662
rect 10600 6598 10652 6604
rect 10508 6384 10560 6390
rect 10508 6326 10560 6332
rect 10508 6248 10560 6254
rect 10428 6196 10508 6202
rect 10428 6190 10560 6196
rect 10428 6174 10548 6190
rect 9588 6112 9640 6118
rect 9588 6054 9640 6060
rect 10428 5914 10456 6174
rect 10612 6118 10640 6598
rect 10704 6322 10732 6870
rect 10888 6798 10916 7534
rect 11060 7482 11112 7488
rect 11164 7342 11192 7890
rect 11244 7744 11296 7750
rect 11244 7686 11296 7692
rect 11256 7478 11284 7686
rect 11244 7472 11296 7478
rect 11244 7414 11296 7420
rect 11152 7336 11204 7342
rect 11152 7278 11204 7284
rect 10784 6792 10836 6798
rect 10784 6734 10836 6740
rect 10876 6792 10928 6798
rect 11164 6746 11192 7278
rect 11244 6996 11296 7002
rect 11244 6938 11296 6944
rect 10876 6734 10928 6740
rect 10796 6390 10824 6734
rect 11072 6718 11192 6746
rect 11072 6662 11100 6718
rect 11060 6656 11112 6662
rect 11060 6598 11112 6604
rect 10784 6384 10836 6390
rect 10784 6326 10836 6332
rect 11072 6322 11100 6598
rect 11256 6458 11284 6938
rect 11348 6730 11376 8502
rect 11624 7954 11652 8978
rect 11716 8906 11744 9998
rect 11808 9926 11836 10134
rect 11900 10130 11928 11070
rect 12072 11018 12124 11024
rect 12348 11076 12400 11082
rect 12348 11018 12400 11024
rect 12256 11008 12308 11014
rect 12256 10950 12308 10956
rect 12268 10470 12296 10950
rect 12360 10470 12388 11018
rect 12532 11008 12584 11014
rect 12532 10950 12584 10956
rect 12544 10742 12572 10950
rect 12638 10908 12946 10917
rect 12638 10906 12644 10908
rect 12700 10906 12724 10908
rect 12780 10906 12804 10908
rect 12860 10906 12884 10908
rect 12940 10906 12946 10908
rect 12700 10854 12702 10906
rect 12882 10854 12884 10906
rect 12638 10852 12644 10854
rect 12700 10852 12724 10854
rect 12780 10852 12804 10854
rect 12860 10852 12884 10854
rect 12940 10852 12946 10854
rect 12638 10843 12946 10852
rect 12532 10736 12584 10742
rect 12532 10678 12584 10684
rect 12256 10464 12308 10470
rect 12256 10406 12308 10412
rect 12348 10464 12400 10470
rect 12348 10406 12400 10412
rect 11978 10364 12286 10373
rect 11978 10362 11984 10364
rect 12040 10362 12064 10364
rect 12120 10362 12144 10364
rect 12200 10362 12224 10364
rect 12280 10362 12286 10364
rect 12040 10310 12042 10362
rect 12222 10310 12224 10362
rect 11978 10308 11984 10310
rect 12040 10308 12064 10310
rect 12120 10308 12144 10310
rect 12200 10308 12224 10310
rect 12280 10308 12286 10310
rect 11978 10299 12286 10308
rect 11888 10124 11940 10130
rect 11888 10066 11940 10072
rect 12072 10056 12124 10062
rect 12072 9998 12124 10004
rect 11796 9920 11848 9926
rect 11796 9862 11848 9868
rect 11888 9920 11940 9926
rect 11888 9862 11940 9868
rect 11704 8900 11756 8906
rect 11704 8842 11756 8848
rect 11612 7948 11664 7954
rect 11612 7890 11664 7896
rect 11624 7410 11652 7890
rect 11716 7886 11744 8842
rect 11704 7880 11756 7886
rect 11704 7822 11756 7828
rect 11716 7546 11744 7822
rect 11808 7818 11836 9862
rect 11900 8566 11928 9862
rect 12084 9722 12112 9998
rect 12360 9926 12388 10406
rect 12532 10124 12584 10130
rect 12532 10066 12584 10072
rect 12544 9994 12572 10066
rect 13268 10056 13320 10062
rect 13268 9998 13320 10004
rect 12532 9988 12584 9994
rect 12532 9930 12584 9936
rect 12348 9920 12400 9926
rect 12348 9862 12400 9868
rect 12638 9820 12946 9829
rect 12638 9818 12644 9820
rect 12700 9818 12724 9820
rect 12780 9818 12804 9820
rect 12860 9818 12884 9820
rect 12940 9818 12946 9820
rect 12700 9766 12702 9818
rect 12882 9766 12884 9818
rect 12638 9764 12644 9766
rect 12700 9764 12724 9766
rect 12780 9764 12804 9766
rect 12860 9764 12884 9766
rect 12940 9764 12946 9766
rect 12638 9755 12946 9764
rect 12072 9716 12124 9722
rect 12072 9658 12124 9664
rect 12348 9648 12400 9654
rect 12348 9590 12400 9596
rect 11978 9276 12286 9285
rect 11978 9274 11984 9276
rect 12040 9274 12064 9276
rect 12120 9274 12144 9276
rect 12200 9274 12224 9276
rect 12280 9274 12286 9276
rect 12040 9222 12042 9274
rect 12222 9222 12224 9274
rect 11978 9220 11984 9222
rect 12040 9220 12064 9222
rect 12120 9220 12144 9222
rect 12200 9220 12224 9222
rect 12280 9220 12286 9222
rect 11978 9211 12286 9220
rect 12360 9178 12388 9590
rect 13280 9518 13308 9998
rect 13268 9512 13320 9518
rect 13268 9454 13320 9460
rect 12348 9172 12400 9178
rect 12348 9114 12400 9120
rect 13280 9042 13308 9454
rect 13268 9036 13320 9042
rect 13268 8978 13320 8984
rect 12348 8968 12400 8974
rect 12348 8910 12400 8916
rect 11888 8560 11940 8566
rect 11888 8502 11940 8508
rect 11978 8188 12286 8197
rect 11978 8186 11984 8188
rect 12040 8186 12064 8188
rect 12120 8186 12144 8188
rect 12200 8186 12224 8188
rect 12280 8186 12286 8188
rect 12040 8134 12042 8186
rect 12222 8134 12224 8186
rect 11978 8132 11984 8134
rect 12040 8132 12064 8134
rect 12120 8132 12144 8134
rect 12200 8132 12224 8134
rect 12280 8132 12286 8134
rect 11978 8123 12286 8132
rect 12360 8022 12388 8910
rect 12638 8732 12946 8741
rect 12638 8730 12644 8732
rect 12700 8730 12724 8732
rect 12780 8730 12804 8732
rect 12860 8730 12884 8732
rect 12940 8730 12946 8732
rect 12700 8678 12702 8730
rect 12882 8678 12884 8730
rect 12638 8676 12644 8678
rect 12700 8676 12724 8678
rect 12780 8676 12804 8678
rect 12860 8676 12884 8678
rect 12940 8676 12946 8678
rect 12638 8667 12946 8676
rect 12348 8016 12400 8022
rect 12348 7958 12400 7964
rect 11796 7812 11848 7818
rect 11796 7754 11848 7760
rect 11704 7540 11756 7546
rect 11704 7482 11756 7488
rect 11808 7410 11836 7754
rect 12256 7744 12308 7750
rect 12256 7686 12308 7692
rect 11428 7404 11480 7410
rect 11428 7346 11480 7352
rect 11612 7404 11664 7410
rect 11612 7346 11664 7352
rect 11796 7404 11848 7410
rect 11796 7346 11848 7352
rect 11440 6798 11468 7346
rect 12268 7206 12296 7686
rect 12360 7460 12388 7958
rect 12638 7644 12946 7653
rect 12638 7642 12644 7644
rect 12700 7642 12724 7644
rect 12780 7642 12804 7644
rect 12860 7642 12884 7644
rect 12940 7642 12946 7644
rect 12700 7590 12702 7642
rect 12882 7590 12884 7642
rect 12638 7588 12644 7590
rect 12700 7588 12724 7590
rect 12780 7588 12804 7590
rect 12860 7588 12884 7590
rect 12940 7588 12946 7590
rect 12638 7579 12946 7588
rect 12532 7472 12584 7478
rect 12360 7432 12532 7460
rect 12532 7414 12584 7420
rect 13268 7336 13320 7342
rect 13268 7278 13320 7284
rect 12256 7200 12308 7206
rect 12256 7142 12308 7148
rect 12532 7200 12584 7206
rect 12532 7142 12584 7148
rect 12900 7200 12952 7206
rect 12900 7142 12952 7148
rect 13176 7200 13228 7206
rect 13176 7142 13228 7148
rect 11978 7100 12286 7109
rect 11978 7098 11984 7100
rect 12040 7098 12064 7100
rect 12120 7098 12144 7100
rect 12200 7098 12224 7100
rect 12280 7098 12286 7100
rect 12040 7046 12042 7098
rect 12222 7046 12224 7098
rect 11978 7044 11984 7046
rect 12040 7044 12064 7046
rect 12120 7044 12144 7046
rect 12200 7044 12224 7046
rect 12280 7044 12286 7046
rect 11978 7035 12286 7044
rect 12544 7002 12572 7142
rect 12532 6996 12584 7002
rect 12532 6938 12584 6944
rect 12912 6798 12940 7142
rect 11428 6792 11480 6798
rect 11428 6734 11480 6740
rect 12900 6792 12952 6798
rect 12900 6734 12952 6740
rect 11336 6724 11388 6730
rect 11336 6666 11388 6672
rect 12638 6556 12946 6565
rect 12638 6554 12644 6556
rect 12700 6554 12724 6556
rect 12780 6554 12804 6556
rect 12860 6554 12884 6556
rect 12940 6554 12946 6556
rect 12700 6502 12702 6554
rect 12882 6502 12884 6554
rect 12638 6500 12644 6502
rect 12700 6500 12724 6502
rect 12780 6500 12804 6502
rect 12860 6500 12884 6502
rect 12940 6500 12946 6502
rect 12638 6491 12946 6500
rect 11244 6452 11296 6458
rect 11244 6394 11296 6400
rect 13188 6390 13216 7142
rect 13280 6866 13308 7278
rect 13268 6860 13320 6866
rect 13268 6802 13320 6808
rect 13176 6384 13228 6390
rect 13176 6326 13228 6332
rect 10692 6316 10744 6322
rect 10692 6258 10744 6264
rect 11060 6316 11112 6322
rect 11060 6258 11112 6264
rect 11796 6248 11848 6254
rect 11796 6190 11848 6196
rect 10600 6112 10652 6118
rect 10600 6054 10652 6060
rect 10784 6112 10836 6118
rect 10784 6054 10836 6060
rect 10416 5908 10468 5914
rect 10416 5850 10468 5856
rect 9487 5468 9795 5477
rect 9487 5466 9493 5468
rect 9549 5466 9573 5468
rect 9629 5466 9653 5468
rect 9709 5466 9733 5468
rect 9789 5466 9795 5468
rect 9549 5414 9551 5466
rect 9731 5414 9733 5466
rect 9487 5412 9493 5414
rect 9549 5412 9573 5414
rect 9629 5412 9653 5414
rect 9709 5412 9733 5414
rect 9789 5412 9795 5414
rect 9487 5403 9795 5412
rect 10428 5386 10456 5850
rect 10796 5710 10824 6054
rect 11808 5914 11836 6190
rect 11978 6012 12286 6021
rect 11978 6010 11984 6012
rect 12040 6010 12064 6012
rect 12120 6010 12144 6012
rect 12200 6010 12224 6012
rect 12280 6010 12286 6012
rect 12040 5958 12042 6010
rect 12222 5958 12224 6010
rect 11978 5956 11984 5958
rect 12040 5956 12064 5958
rect 12120 5956 12144 5958
rect 12200 5956 12224 5958
rect 12280 5956 12286 5958
rect 11978 5947 12286 5956
rect 11796 5908 11848 5914
rect 11796 5850 11848 5856
rect 10784 5704 10836 5710
rect 10784 5646 10836 5652
rect 12638 5468 12946 5477
rect 12638 5466 12644 5468
rect 12700 5466 12724 5468
rect 12780 5466 12804 5468
rect 12860 5466 12884 5468
rect 12940 5466 12946 5468
rect 12700 5414 12702 5466
rect 12882 5414 12884 5466
rect 12638 5412 12644 5414
rect 12700 5412 12724 5414
rect 12780 5412 12804 5414
rect 12860 5412 12884 5414
rect 12940 5412 12946 5414
rect 12638 5403 12946 5412
rect 10336 5358 10456 5386
rect 9680 5024 9732 5030
rect 9680 4966 9732 4972
rect 9692 4622 9720 4966
rect 10336 4690 10364 5358
rect 10784 5024 10836 5030
rect 10784 4966 10836 4972
rect 9956 4684 10008 4690
rect 9956 4626 10008 4632
rect 10324 4684 10376 4690
rect 10324 4626 10376 4632
rect 9220 4616 9272 4622
rect 9220 4558 9272 4564
rect 9312 4616 9364 4622
rect 9312 4558 9364 4564
rect 9680 4616 9732 4622
rect 9680 4558 9732 4564
rect 8668 4480 8720 4486
rect 8668 4422 8720 4428
rect 9128 4480 9180 4486
rect 9128 4422 9180 4428
rect 8484 3596 8536 3602
rect 8484 3538 8536 3544
rect 8392 3188 8444 3194
rect 8392 3130 8444 3136
rect 8496 3126 8524 3538
rect 8576 3528 8628 3534
rect 8576 3470 8628 3476
rect 8484 3120 8536 3126
rect 8484 3062 8536 3068
rect 8588 3058 8616 3470
rect 8680 3194 8708 4422
rect 9140 4078 9168 4422
rect 9128 4072 9180 4078
rect 9128 4014 9180 4020
rect 8827 3836 9135 3845
rect 8827 3834 8833 3836
rect 8889 3834 8913 3836
rect 8969 3834 8993 3836
rect 9049 3834 9073 3836
rect 9129 3834 9135 3836
rect 8889 3782 8891 3834
rect 9071 3782 9073 3834
rect 8827 3780 8833 3782
rect 8889 3780 8913 3782
rect 8969 3780 8993 3782
rect 9049 3780 9073 3782
rect 9129 3780 9135 3782
rect 8827 3771 9135 3780
rect 9232 3194 9260 4558
rect 9312 4480 9364 4486
rect 9312 4422 9364 4428
rect 8668 3188 8720 3194
rect 8668 3130 8720 3136
rect 9220 3188 9272 3194
rect 9220 3130 9272 3136
rect 7932 3052 7984 3058
rect 7932 2994 7984 3000
rect 8576 3052 8628 3058
rect 8576 2994 8628 3000
rect 9324 2854 9352 4422
rect 9487 4380 9795 4389
rect 9487 4378 9493 4380
rect 9549 4378 9573 4380
rect 9629 4378 9653 4380
rect 9709 4378 9733 4380
rect 9789 4378 9795 4380
rect 9549 4326 9551 4378
rect 9731 4326 9733 4378
rect 9487 4324 9493 4326
rect 9549 4324 9573 4326
rect 9629 4324 9653 4326
rect 9709 4324 9733 4326
rect 9789 4324 9795 4326
rect 9487 4315 9795 4324
rect 9968 4282 9996 4626
rect 10048 4616 10100 4622
rect 10048 4558 10100 4564
rect 9956 4276 10008 4282
rect 9956 4218 10008 4224
rect 9772 4140 9824 4146
rect 9772 4082 9824 4088
rect 9404 3936 9456 3942
rect 9404 3878 9456 3884
rect 9416 3194 9444 3878
rect 9784 3602 9812 4082
rect 9968 3942 9996 4218
rect 9956 3936 10008 3942
rect 9956 3878 10008 3884
rect 9772 3596 9824 3602
rect 9772 3538 9824 3544
rect 9487 3292 9795 3301
rect 9487 3290 9493 3292
rect 9549 3290 9573 3292
rect 9629 3290 9653 3292
rect 9709 3290 9733 3292
rect 9789 3290 9795 3292
rect 9549 3238 9551 3290
rect 9731 3238 9733 3290
rect 9487 3236 9493 3238
rect 9549 3236 9573 3238
rect 9629 3236 9653 3238
rect 9709 3236 9733 3238
rect 9789 3236 9795 3238
rect 9487 3227 9795 3236
rect 10060 3194 10088 4558
rect 10140 4548 10192 4554
rect 10140 4490 10192 4496
rect 10152 4078 10180 4490
rect 10336 4214 10364 4626
rect 10796 4486 10824 4966
rect 11978 4924 12286 4933
rect 11978 4922 11984 4924
rect 12040 4922 12064 4924
rect 12120 4922 12144 4924
rect 12200 4922 12224 4924
rect 12280 4922 12286 4924
rect 12040 4870 12042 4922
rect 12222 4870 12224 4922
rect 11978 4868 11984 4870
rect 12040 4868 12064 4870
rect 12120 4868 12144 4870
rect 12200 4868 12224 4870
rect 12280 4868 12286 4870
rect 11978 4859 12286 4868
rect 10968 4684 11020 4690
rect 10968 4626 11020 4632
rect 10784 4480 10836 4486
rect 10784 4422 10836 4428
rect 10692 4276 10744 4282
rect 10692 4218 10744 4224
rect 10324 4208 10376 4214
rect 10324 4150 10376 4156
rect 10416 4208 10468 4214
rect 10416 4150 10468 4156
rect 10140 4072 10192 4078
rect 10428 4060 10456 4150
rect 10192 4032 10456 4060
rect 10140 4014 10192 4020
rect 9404 3188 9456 3194
rect 9404 3130 9456 3136
rect 10048 3188 10100 3194
rect 10048 3130 10100 3136
rect 9416 2922 9444 3130
rect 9404 2916 9456 2922
rect 9404 2858 9456 2864
rect 9312 2848 9364 2854
rect 9312 2790 9364 2796
rect 8827 2748 9135 2757
rect 8827 2746 8833 2748
rect 8889 2746 8913 2748
rect 8969 2746 8993 2748
rect 9049 2746 9073 2748
rect 9129 2746 9135 2748
rect 8889 2694 8891 2746
rect 9071 2694 9073 2746
rect 8827 2692 8833 2694
rect 8889 2692 8913 2694
rect 8969 2692 8993 2694
rect 9049 2692 9073 2694
rect 9129 2692 9135 2694
rect 8827 2683 9135 2692
rect 4160 2644 4212 2650
rect 4160 2586 4212 2592
rect 7380 2644 7432 2650
rect 7380 2586 7432 2592
rect 10152 2514 10180 4014
rect 10704 3738 10732 4218
rect 10796 4146 10824 4422
rect 10980 4282 11008 4626
rect 12992 4616 13044 4622
rect 12992 4558 13044 4564
rect 13176 4616 13228 4622
rect 13176 4558 13228 4564
rect 12440 4480 12492 4486
rect 12440 4422 12492 4428
rect 10968 4276 11020 4282
rect 10968 4218 11020 4224
rect 10784 4140 10836 4146
rect 10784 4082 10836 4088
rect 11152 4140 11204 4146
rect 11152 4082 11204 4088
rect 10692 3732 10744 3738
rect 10692 3674 10744 3680
rect 10704 2990 10732 3674
rect 10232 2984 10284 2990
rect 10232 2926 10284 2932
rect 10692 2984 10744 2990
rect 10692 2926 10744 2932
rect 10140 2508 10192 2514
rect 10140 2450 10192 2456
rect 10244 2446 10272 2926
rect 10796 2446 10824 4082
rect 11164 3942 11192 4082
rect 11152 3936 11204 3942
rect 11152 3878 11204 3884
rect 11520 3936 11572 3942
rect 11520 3878 11572 3884
rect 11164 3058 11192 3878
rect 11532 3602 11560 3878
rect 11978 3836 12286 3845
rect 11978 3834 11984 3836
rect 12040 3834 12064 3836
rect 12120 3834 12144 3836
rect 12200 3834 12224 3836
rect 12280 3834 12286 3836
rect 12040 3782 12042 3834
rect 12222 3782 12224 3834
rect 11978 3780 11984 3782
rect 12040 3780 12064 3782
rect 12120 3780 12144 3782
rect 12200 3780 12224 3782
rect 12280 3780 12286 3782
rect 11978 3771 12286 3780
rect 11520 3596 11572 3602
rect 11520 3538 11572 3544
rect 12452 3466 12480 4422
rect 12638 4380 12946 4389
rect 12638 4378 12644 4380
rect 12700 4378 12724 4380
rect 12780 4378 12804 4380
rect 12860 4378 12884 4380
rect 12940 4378 12946 4380
rect 12700 4326 12702 4378
rect 12882 4326 12884 4378
rect 12638 4324 12644 4326
rect 12700 4324 12724 4326
rect 12780 4324 12804 4326
rect 12860 4324 12884 4326
rect 12940 4324 12946 4326
rect 12638 4315 12946 4324
rect 13004 4146 13032 4558
rect 13084 4480 13136 4486
rect 13084 4422 13136 4428
rect 13096 4146 13124 4422
rect 12992 4140 13044 4146
rect 12992 4082 13044 4088
rect 13084 4140 13136 4146
rect 13084 4082 13136 4088
rect 13188 4078 13216 4558
rect 13268 4480 13320 4486
rect 13268 4422 13320 4428
rect 13280 4185 13308 4422
rect 13266 4176 13322 4185
rect 13266 4111 13322 4120
rect 13176 4072 13228 4078
rect 13176 4014 13228 4020
rect 12532 4004 12584 4010
rect 12532 3946 12584 3952
rect 12544 3738 12572 3946
rect 12532 3732 12584 3738
rect 12532 3674 12584 3680
rect 13360 3528 13412 3534
rect 13358 3496 13360 3505
rect 13412 3496 13414 3505
rect 12440 3460 12492 3466
rect 13358 3431 13414 3440
rect 12440 3402 12492 3408
rect 12638 3292 12946 3301
rect 12638 3290 12644 3292
rect 12700 3290 12724 3292
rect 12780 3290 12804 3292
rect 12860 3290 12884 3292
rect 12940 3290 12946 3292
rect 12700 3238 12702 3290
rect 12882 3238 12884 3290
rect 12638 3236 12644 3238
rect 12700 3236 12724 3238
rect 12780 3236 12804 3238
rect 12860 3236 12884 3238
rect 12940 3236 12946 3238
rect 12638 3227 12946 3236
rect 11152 3052 11204 3058
rect 11152 2994 11204 3000
rect 13360 2984 13412 2990
rect 13360 2926 13412 2932
rect 13372 2825 13400 2926
rect 13358 2816 13414 2825
rect 11978 2748 12286 2757
rect 13358 2751 13414 2760
rect 11978 2746 11984 2748
rect 12040 2746 12064 2748
rect 12120 2746 12144 2748
rect 12200 2746 12224 2748
rect 12280 2746 12286 2748
rect 12040 2694 12042 2746
rect 12222 2694 12224 2746
rect 11978 2692 11984 2694
rect 12040 2692 12064 2694
rect 12120 2692 12144 2694
rect 12200 2692 12224 2694
rect 12280 2692 12286 2694
rect 11978 2683 12286 2692
rect 3608 2440 3660 2446
rect 3608 2382 3660 2388
rect 7104 2440 7156 2446
rect 7104 2382 7156 2388
rect 10232 2440 10284 2446
rect 10232 2382 10284 2388
rect 10784 2440 10836 2446
rect 10784 2382 10836 2388
rect 3185 2204 3493 2213
rect 3185 2202 3191 2204
rect 3247 2202 3271 2204
rect 3327 2202 3351 2204
rect 3407 2202 3431 2204
rect 3487 2202 3493 2204
rect 3247 2150 3249 2202
rect 3429 2150 3431 2202
rect 3185 2148 3191 2150
rect 3247 2148 3271 2150
rect 3327 2148 3351 2150
rect 3407 2148 3431 2150
rect 3487 2148 3493 2150
rect 3185 2139 3493 2148
rect 6336 2204 6644 2213
rect 6336 2202 6342 2204
rect 6398 2202 6422 2204
rect 6478 2202 6502 2204
rect 6558 2202 6582 2204
rect 6638 2202 6644 2204
rect 6398 2150 6400 2202
rect 6580 2150 6582 2202
rect 6336 2148 6342 2150
rect 6398 2148 6422 2150
rect 6478 2148 6502 2150
rect 6558 2148 6582 2150
rect 6638 2148 6644 2150
rect 6336 2139 6644 2148
rect 7116 800 7144 2382
rect 9036 2304 9088 2310
rect 9036 2246 9088 2252
rect 9864 2304 9916 2310
rect 9864 2246 9916 2252
rect 10324 2304 10376 2310
rect 10324 2246 10376 2252
rect 9048 800 9076 2246
rect 9487 2204 9795 2213
rect 9487 2202 9493 2204
rect 9549 2202 9573 2204
rect 9629 2202 9653 2204
rect 9709 2202 9733 2204
rect 9789 2202 9795 2204
rect 9549 2150 9551 2202
rect 9731 2150 9733 2202
rect 9487 2148 9493 2150
rect 9549 2148 9573 2150
rect 9629 2148 9653 2150
rect 9709 2148 9733 2150
rect 9789 2148 9795 2150
rect 9487 2139 9795 2148
rect 9876 1170 9904 2246
rect 9692 1142 9904 1170
rect 9692 800 9720 1142
rect 10336 800 10364 2246
rect 12638 2204 12946 2213
rect 12638 2202 12644 2204
rect 12700 2202 12724 2204
rect 12780 2202 12804 2204
rect 12860 2202 12884 2204
rect 12940 2202 12946 2204
rect 12700 2150 12702 2202
rect 12882 2150 12884 2202
rect 12638 2148 12644 2150
rect 12700 2148 12724 2150
rect 12780 2148 12804 2150
rect 12860 2148 12884 2150
rect 12940 2148 12946 2150
rect 12638 2139 12946 2148
rect 7102 0 7158 800
rect 9034 0 9090 800
rect 9678 0 9734 800
rect 10322 0 10378 800
<< via2 >>
rect 2531 14714 2587 14716
rect 2611 14714 2667 14716
rect 2691 14714 2747 14716
rect 2771 14714 2827 14716
rect 2531 14662 2577 14714
rect 2577 14662 2587 14714
rect 2611 14662 2641 14714
rect 2641 14662 2653 14714
rect 2653 14662 2667 14714
rect 2691 14662 2705 14714
rect 2705 14662 2717 14714
rect 2717 14662 2747 14714
rect 2771 14662 2781 14714
rect 2781 14662 2827 14714
rect 2531 14660 2587 14662
rect 2611 14660 2667 14662
rect 2691 14660 2747 14662
rect 2771 14660 2827 14662
rect 5682 14714 5738 14716
rect 5762 14714 5818 14716
rect 5842 14714 5898 14716
rect 5922 14714 5978 14716
rect 5682 14662 5728 14714
rect 5728 14662 5738 14714
rect 5762 14662 5792 14714
rect 5792 14662 5804 14714
rect 5804 14662 5818 14714
rect 5842 14662 5856 14714
rect 5856 14662 5868 14714
rect 5868 14662 5898 14714
rect 5922 14662 5932 14714
rect 5932 14662 5978 14714
rect 5682 14660 5738 14662
rect 5762 14660 5818 14662
rect 5842 14660 5898 14662
rect 5922 14660 5978 14662
rect 8833 14714 8889 14716
rect 8913 14714 8969 14716
rect 8993 14714 9049 14716
rect 9073 14714 9129 14716
rect 8833 14662 8879 14714
rect 8879 14662 8889 14714
rect 8913 14662 8943 14714
rect 8943 14662 8955 14714
rect 8955 14662 8969 14714
rect 8993 14662 9007 14714
rect 9007 14662 9019 14714
rect 9019 14662 9049 14714
rect 9073 14662 9083 14714
rect 9083 14662 9129 14714
rect 8833 14660 8889 14662
rect 8913 14660 8969 14662
rect 8993 14660 9049 14662
rect 9073 14660 9129 14662
rect 11984 14714 12040 14716
rect 12064 14714 12120 14716
rect 12144 14714 12200 14716
rect 12224 14714 12280 14716
rect 11984 14662 12030 14714
rect 12030 14662 12040 14714
rect 12064 14662 12094 14714
rect 12094 14662 12106 14714
rect 12106 14662 12120 14714
rect 12144 14662 12158 14714
rect 12158 14662 12170 14714
rect 12170 14662 12200 14714
rect 12224 14662 12234 14714
rect 12234 14662 12280 14714
rect 11984 14660 12040 14662
rect 12064 14660 12120 14662
rect 12144 14660 12200 14662
rect 12224 14660 12280 14662
rect 3191 14170 3247 14172
rect 3271 14170 3327 14172
rect 3351 14170 3407 14172
rect 3431 14170 3487 14172
rect 3191 14118 3237 14170
rect 3237 14118 3247 14170
rect 3271 14118 3301 14170
rect 3301 14118 3313 14170
rect 3313 14118 3327 14170
rect 3351 14118 3365 14170
rect 3365 14118 3377 14170
rect 3377 14118 3407 14170
rect 3431 14118 3441 14170
rect 3441 14118 3487 14170
rect 3191 14116 3247 14118
rect 3271 14116 3327 14118
rect 3351 14116 3407 14118
rect 3431 14116 3487 14118
rect 6342 14170 6398 14172
rect 6422 14170 6478 14172
rect 6502 14170 6558 14172
rect 6582 14170 6638 14172
rect 6342 14118 6388 14170
rect 6388 14118 6398 14170
rect 6422 14118 6452 14170
rect 6452 14118 6464 14170
rect 6464 14118 6478 14170
rect 6502 14118 6516 14170
rect 6516 14118 6528 14170
rect 6528 14118 6558 14170
rect 6582 14118 6592 14170
rect 6592 14118 6638 14170
rect 6342 14116 6398 14118
rect 6422 14116 6478 14118
rect 6502 14116 6558 14118
rect 6582 14116 6638 14118
rect 9493 14170 9549 14172
rect 9573 14170 9629 14172
rect 9653 14170 9709 14172
rect 9733 14170 9789 14172
rect 9493 14118 9539 14170
rect 9539 14118 9549 14170
rect 9573 14118 9603 14170
rect 9603 14118 9615 14170
rect 9615 14118 9629 14170
rect 9653 14118 9667 14170
rect 9667 14118 9679 14170
rect 9679 14118 9709 14170
rect 9733 14118 9743 14170
rect 9743 14118 9789 14170
rect 9493 14116 9549 14118
rect 9573 14116 9629 14118
rect 9653 14116 9709 14118
rect 9733 14116 9789 14118
rect 12644 14170 12700 14172
rect 12724 14170 12780 14172
rect 12804 14170 12860 14172
rect 12884 14170 12940 14172
rect 12644 14118 12690 14170
rect 12690 14118 12700 14170
rect 12724 14118 12754 14170
rect 12754 14118 12766 14170
rect 12766 14118 12780 14170
rect 12804 14118 12818 14170
rect 12818 14118 12830 14170
rect 12830 14118 12860 14170
rect 12884 14118 12894 14170
rect 12894 14118 12940 14170
rect 12644 14116 12700 14118
rect 12724 14116 12780 14118
rect 12804 14116 12860 14118
rect 12884 14116 12940 14118
rect 1398 13640 1454 13696
rect 2531 13626 2587 13628
rect 2611 13626 2667 13628
rect 2691 13626 2747 13628
rect 2771 13626 2827 13628
rect 2531 13574 2577 13626
rect 2577 13574 2587 13626
rect 2611 13574 2641 13626
rect 2641 13574 2653 13626
rect 2653 13574 2667 13626
rect 2691 13574 2705 13626
rect 2705 13574 2717 13626
rect 2717 13574 2747 13626
rect 2771 13574 2781 13626
rect 2781 13574 2827 13626
rect 2531 13572 2587 13574
rect 2611 13572 2667 13574
rect 2691 13572 2747 13574
rect 2771 13572 2827 13574
rect 846 13132 848 13152
rect 848 13132 900 13152
rect 900 13132 902 13152
rect 846 13096 902 13132
rect 3191 13082 3247 13084
rect 3271 13082 3327 13084
rect 3351 13082 3407 13084
rect 3431 13082 3487 13084
rect 3191 13030 3237 13082
rect 3237 13030 3247 13082
rect 3271 13030 3301 13082
rect 3301 13030 3313 13082
rect 3313 13030 3327 13082
rect 3351 13030 3365 13082
rect 3365 13030 3377 13082
rect 3377 13030 3407 13082
rect 3431 13030 3441 13082
rect 3441 13030 3487 13082
rect 3191 13028 3247 13030
rect 3271 13028 3327 13030
rect 3351 13028 3407 13030
rect 3431 13028 3487 13030
rect 2531 12538 2587 12540
rect 2611 12538 2667 12540
rect 2691 12538 2747 12540
rect 2771 12538 2827 12540
rect 2531 12486 2577 12538
rect 2577 12486 2587 12538
rect 2611 12486 2641 12538
rect 2641 12486 2653 12538
rect 2653 12486 2667 12538
rect 2691 12486 2705 12538
rect 2705 12486 2717 12538
rect 2717 12486 2747 12538
rect 2771 12486 2781 12538
rect 2781 12486 2827 12538
rect 2531 12484 2587 12486
rect 2611 12484 2667 12486
rect 2691 12484 2747 12486
rect 2771 12484 2827 12486
rect 3191 11994 3247 11996
rect 3271 11994 3327 11996
rect 3351 11994 3407 11996
rect 3431 11994 3487 11996
rect 3191 11942 3237 11994
rect 3237 11942 3247 11994
rect 3271 11942 3301 11994
rect 3301 11942 3313 11994
rect 3313 11942 3327 11994
rect 3351 11942 3365 11994
rect 3365 11942 3377 11994
rect 3377 11942 3407 11994
rect 3431 11942 3441 11994
rect 3441 11942 3487 11994
rect 3191 11940 3247 11942
rect 3271 11940 3327 11942
rect 3351 11940 3407 11942
rect 3431 11940 3487 11942
rect 2531 11450 2587 11452
rect 2611 11450 2667 11452
rect 2691 11450 2747 11452
rect 2771 11450 2827 11452
rect 2531 11398 2577 11450
rect 2577 11398 2587 11450
rect 2611 11398 2641 11450
rect 2641 11398 2653 11450
rect 2653 11398 2667 11450
rect 2691 11398 2705 11450
rect 2705 11398 2717 11450
rect 2717 11398 2747 11450
rect 2771 11398 2781 11450
rect 2781 11398 2827 11450
rect 2531 11396 2587 11398
rect 2611 11396 2667 11398
rect 2691 11396 2747 11398
rect 2771 11396 2827 11398
rect 2531 10362 2587 10364
rect 2611 10362 2667 10364
rect 2691 10362 2747 10364
rect 2771 10362 2827 10364
rect 2531 10310 2577 10362
rect 2577 10310 2587 10362
rect 2611 10310 2641 10362
rect 2641 10310 2653 10362
rect 2653 10310 2667 10362
rect 2691 10310 2705 10362
rect 2705 10310 2717 10362
rect 2717 10310 2747 10362
rect 2771 10310 2781 10362
rect 2781 10310 2827 10362
rect 2531 10308 2587 10310
rect 2611 10308 2667 10310
rect 2691 10308 2747 10310
rect 2771 10308 2827 10310
rect 3191 10906 3247 10908
rect 3271 10906 3327 10908
rect 3351 10906 3407 10908
rect 3431 10906 3487 10908
rect 3191 10854 3237 10906
rect 3237 10854 3247 10906
rect 3271 10854 3301 10906
rect 3301 10854 3313 10906
rect 3313 10854 3327 10906
rect 3351 10854 3365 10906
rect 3365 10854 3377 10906
rect 3377 10854 3407 10906
rect 3431 10854 3441 10906
rect 3441 10854 3487 10906
rect 3191 10852 3247 10854
rect 3271 10852 3327 10854
rect 3351 10852 3407 10854
rect 3431 10852 3487 10854
rect 2531 9274 2587 9276
rect 2611 9274 2667 9276
rect 2691 9274 2747 9276
rect 2771 9274 2827 9276
rect 2531 9222 2577 9274
rect 2577 9222 2587 9274
rect 2611 9222 2641 9274
rect 2641 9222 2653 9274
rect 2653 9222 2667 9274
rect 2691 9222 2705 9274
rect 2705 9222 2717 9274
rect 2717 9222 2747 9274
rect 2771 9222 2781 9274
rect 2781 9222 2827 9274
rect 2531 9220 2587 9222
rect 2611 9220 2667 9222
rect 2691 9220 2747 9222
rect 2771 9220 2827 9222
rect 2531 8186 2587 8188
rect 2611 8186 2667 8188
rect 2691 8186 2747 8188
rect 2771 8186 2827 8188
rect 2531 8134 2577 8186
rect 2577 8134 2587 8186
rect 2611 8134 2641 8186
rect 2641 8134 2653 8186
rect 2653 8134 2667 8186
rect 2691 8134 2705 8186
rect 2705 8134 2717 8186
rect 2717 8134 2747 8186
rect 2771 8134 2781 8186
rect 2781 8134 2827 8186
rect 2531 8132 2587 8134
rect 2611 8132 2667 8134
rect 2691 8132 2747 8134
rect 2771 8132 2827 8134
rect 3191 9818 3247 9820
rect 3271 9818 3327 9820
rect 3351 9818 3407 9820
rect 3431 9818 3487 9820
rect 3191 9766 3237 9818
rect 3237 9766 3247 9818
rect 3271 9766 3301 9818
rect 3301 9766 3313 9818
rect 3313 9766 3327 9818
rect 3351 9766 3365 9818
rect 3365 9766 3377 9818
rect 3377 9766 3407 9818
rect 3431 9766 3441 9818
rect 3441 9766 3487 9818
rect 3191 9764 3247 9766
rect 3271 9764 3327 9766
rect 3351 9764 3407 9766
rect 3431 9764 3487 9766
rect 5682 13626 5738 13628
rect 5762 13626 5818 13628
rect 5842 13626 5898 13628
rect 5922 13626 5978 13628
rect 5682 13574 5728 13626
rect 5728 13574 5738 13626
rect 5762 13574 5792 13626
rect 5792 13574 5804 13626
rect 5804 13574 5818 13626
rect 5842 13574 5856 13626
rect 5856 13574 5868 13626
rect 5868 13574 5898 13626
rect 5922 13574 5932 13626
rect 5932 13574 5978 13626
rect 5682 13572 5738 13574
rect 5762 13572 5818 13574
rect 5842 13572 5898 13574
rect 5922 13572 5978 13574
rect 5682 12538 5738 12540
rect 5762 12538 5818 12540
rect 5842 12538 5898 12540
rect 5922 12538 5978 12540
rect 5682 12486 5728 12538
rect 5728 12486 5738 12538
rect 5762 12486 5792 12538
rect 5792 12486 5804 12538
rect 5804 12486 5818 12538
rect 5842 12486 5856 12538
rect 5856 12486 5868 12538
rect 5868 12486 5898 12538
rect 5922 12486 5932 12538
rect 5932 12486 5978 12538
rect 5682 12484 5738 12486
rect 5762 12484 5818 12486
rect 5842 12484 5898 12486
rect 5922 12484 5978 12486
rect 6342 13082 6398 13084
rect 6422 13082 6478 13084
rect 6502 13082 6558 13084
rect 6582 13082 6638 13084
rect 6342 13030 6388 13082
rect 6388 13030 6398 13082
rect 6422 13030 6452 13082
rect 6452 13030 6464 13082
rect 6464 13030 6478 13082
rect 6502 13030 6516 13082
rect 6516 13030 6528 13082
rect 6528 13030 6558 13082
rect 6582 13030 6592 13082
rect 6592 13030 6638 13082
rect 6342 13028 6398 13030
rect 6422 13028 6478 13030
rect 6502 13028 6558 13030
rect 6582 13028 6638 13030
rect 6342 11994 6398 11996
rect 6422 11994 6478 11996
rect 6502 11994 6558 11996
rect 6582 11994 6638 11996
rect 6342 11942 6388 11994
rect 6388 11942 6398 11994
rect 6422 11942 6452 11994
rect 6452 11942 6464 11994
rect 6464 11942 6478 11994
rect 6502 11942 6516 11994
rect 6516 11942 6528 11994
rect 6528 11942 6558 11994
rect 6582 11942 6592 11994
rect 6592 11942 6638 11994
rect 6342 11940 6398 11942
rect 6422 11940 6478 11942
rect 6502 11940 6558 11942
rect 6582 11940 6638 11942
rect 5682 11450 5738 11452
rect 5762 11450 5818 11452
rect 5842 11450 5898 11452
rect 5922 11450 5978 11452
rect 5682 11398 5728 11450
rect 5728 11398 5738 11450
rect 5762 11398 5792 11450
rect 5792 11398 5804 11450
rect 5804 11398 5818 11450
rect 5842 11398 5856 11450
rect 5856 11398 5868 11450
rect 5868 11398 5898 11450
rect 5922 11398 5932 11450
rect 5932 11398 5978 11450
rect 5682 11396 5738 11398
rect 5762 11396 5818 11398
rect 5842 11396 5898 11398
rect 5922 11396 5978 11398
rect 6342 10906 6398 10908
rect 6422 10906 6478 10908
rect 6502 10906 6558 10908
rect 6582 10906 6638 10908
rect 6342 10854 6388 10906
rect 6388 10854 6398 10906
rect 6422 10854 6452 10906
rect 6452 10854 6464 10906
rect 6464 10854 6478 10906
rect 6502 10854 6516 10906
rect 6516 10854 6528 10906
rect 6528 10854 6558 10906
rect 6582 10854 6592 10906
rect 6592 10854 6638 10906
rect 6342 10852 6398 10854
rect 6422 10852 6478 10854
rect 6502 10852 6558 10854
rect 6582 10852 6638 10854
rect 8833 13626 8889 13628
rect 8913 13626 8969 13628
rect 8993 13626 9049 13628
rect 9073 13626 9129 13628
rect 8833 13574 8879 13626
rect 8879 13574 8889 13626
rect 8913 13574 8943 13626
rect 8943 13574 8955 13626
rect 8955 13574 8969 13626
rect 8993 13574 9007 13626
rect 9007 13574 9019 13626
rect 9019 13574 9049 13626
rect 9073 13574 9083 13626
rect 9083 13574 9129 13626
rect 8833 13572 8889 13574
rect 8913 13572 8969 13574
rect 8993 13572 9049 13574
rect 9073 13572 9129 13574
rect 5682 10362 5738 10364
rect 5762 10362 5818 10364
rect 5842 10362 5898 10364
rect 5922 10362 5978 10364
rect 5682 10310 5728 10362
rect 5728 10310 5738 10362
rect 5762 10310 5792 10362
rect 5792 10310 5804 10362
rect 5804 10310 5818 10362
rect 5842 10310 5856 10362
rect 5856 10310 5868 10362
rect 5868 10310 5898 10362
rect 5922 10310 5932 10362
rect 5932 10310 5978 10362
rect 5682 10308 5738 10310
rect 5762 10308 5818 10310
rect 5842 10308 5898 10310
rect 5922 10308 5978 10310
rect 6342 9818 6398 9820
rect 6422 9818 6478 9820
rect 6502 9818 6558 9820
rect 6582 9818 6638 9820
rect 6342 9766 6388 9818
rect 6388 9766 6398 9818
rect 6422 9766 6452 9818
rect 6452 9766 6464 9818
rect 6464 9766 6478 9818
rect 6502 9766 6516 9818
rect 6516 9766 6528 9818
rect 6528 9766 6558 9818
rect 6582 9766 6592 9818
rect 6592 9766 6638 9818
rect 6342 9764 6398 9766
rect 6422 9764 6478 9766
rect 6502 9764 6558 9766
rect 6582 9764 6638 9766
rect 6550 9560 6606 9616
rect 3191 8730 3247 8732
rect 3271 8730 3327 8732
rect 3351 8730 3407 8732
rect 3431 8730 3487 8732
rect 3191 8678 3237 8730
rect 3237 8678 3247 8730
rect 3271 8678 3301 8730
rect 3301 8678 3313 8730
rect 3313 8678 3327 8730
rect 3351 8678 3365 8730
rect 3365 8678 3377 8730
rect 3377 8678 3407 8730
rect 3431 8678 3441 8730
rect 3441 8678 3487 8730
rect 3191 8676 3247 8678
rect 3271 8676 3327 8678
rect 3351 8676 3407 8678
rect 3431 8676 3487 8678
rect 2531 7098 2587 7100
rect 2611 7098 2667 7100
rect 2691 7098 2747 7100
rect 2771 7098 2827 7100
rect 2531 7046 2577 7098
rect 2577 7046 2587 7098
rect 2611 7046 2641 7098
rect 2641 7046 2653 7098
rect 2653 7046 2667 7098
rect 2691 7046 2705 7098
rect 2705 7046 2717 7098
rect 2717 7046 2747 7098
rect 2771 7046 2781 7098
rect 2781 7046 2827 7098
rect 2531 7044 2587 7046
rect 2611 7044 2667 7046
rect 2691 7044 2747 7046
rect 2771 7044 2827 7046
rect 2531 6010 2587 6012
rect 2611 6010 2667 6012
rect 2691 6010 2747 6012
rect 2771 6010 2827 6012
rect 2531 5958 2577 6010
rect 2577 5958 2587 6010
rect 2611 5958 2641 6010
rect 2641 5958 2653 6010
rect 2653 5958 2667 6010
rect 2691 5958 2705 6010
rect 2705 5958 2717 6010
rect 2717 5958 2747 6010
rect 2771 5958 2781 6010
rect 2781 5958 2827 6010
rect 2531 5956 2587 5958
rect 2611 5956 2667 5958
rect 2691 5956 2747 5958
rect 2771 5956 2827 5958
rect 3191 7642 3247 7644
rect 3271 7642 3327 7644
rect 3351 7642 3407 7644
rect 3431 7642 3487 7644
rect 3191 7590 3237 7642
rect 3237 7590 3247 7642
rect 3271 7590 3301 7642
rect 3301 7590 3313 7642
rect 3313 7590 3327 7642
rect 3351 7590 3365 7642
rect 3365 7590 3377 7642
rect 3377 7590 3407 7642
rect 3431 7590 3441 7642
rect 3441 7590 3487 7642
rect 3191 7588 3247 7590
rect 3271 7588 3327 7590
rect 3351 7588 3407 7590
rect 3431 7588 3487 7590
rect 3191 6554 3247 6556
rect 3271 6554 3327 6556
rect 3351 6554 3407 6556
rect 3431 6554 3487 6556
rect 3191 6502 3237 6554
rect 3237 6502 3247 6554
rect 3271 6502 3301 6554
rect 3301 6502 3313 6554
rect 3313 6502 3327 6554
rect 3351 6502 3365 6554
rect 3365 6502 3377 6554
rect 3377 6502 3407 6554
rect 3431 6502 3441 6554
rect 3441 6502 3487 6554
rect 3191 6500 3247 6502
rect 3271 6500 3327 6502
rect 3351 6500 3407 6502
rect 3431 6500 3487 6502
rect 5682 9274 5738 9276
rect 5762 9274 5818 9276
rect 5842 9274 5898 9276
rect 5922 9274 5978 9276
rect 5682 9222 5728 9274
rect 5728 9222 5738 9274
rect 5762 9222 5792 9274
rect 5792 9222 5804 9274
rect 5804 9222 5818 9274
rect 5842 9222 5856 9274
rect 5856 9222 5868 9274
rect 5868 9222 5898 9274
rect 5922 9222 5932 9274
rect 5932 9222 5978 9274
rect 5682 9220 5738 9222
rect 5762 9220 5818 9222
rect 5842 9220 5898 9222
rect 5922 9220 5978 9222
rect 6342 8730 6398 8732
rect 6422 8730 6478 8732
rect 6502 8730 6558 8732
rect 6582 8730 6638 8732
rect 6342 8678 6388 8730
rect 6388 8678 6398 8730
rect 6422 8678 6452 8730
rect 6452 8678 6464 8730
rect 6464 8678 6478 8730
rect 6502 8678 6516 8730
rect 6516 8678 6528 8730
rect 6528 8678 6558 8730
rect 6582 8678 6592 8730
rect 6592 8678 6638 8730
rect 6342 8676 6398 8678
rect 6422 8676 6478 8678
rect 6502 8676 6558 8678
rect 6582 8676 6638 8678
rect 5682 8186 5738 8188
rect 5762 8186 5818 8188
rect 5842 8186 5898 8188
rect 5922 8186 5978 8188
rect 5682 8134 5728 8186
rect 5728 8134 5738 8186
rect 5762 8134 5792 8186
rect 5792 8134 5804 8186
rect 5804 8134 5818 8186
rect 5842 8134 5856 8186
rect 5856 8134 5868 8186
rect 5868 8134 5898 8186
rect 5922 8134 5932 8186
rect 5932 8134 5978 8186
rect 5682 8132 5738 8134
rect 5762 8132 5818 8134
rect 5842 8132 5898 8134
rect 5922 8132 5978 8134
rect 6342 7642 6398 7644
rect 6422 7642 6478 7644
rect 6502 7642 6558 7644
rect 6582 7642 6638 7644
rect 6342 7590 6388 7642
rect 6388 7590 6398 7642
rect 6422 7590 6452 7642
rect 6452 7590 6464 7642
rect 6464 7590 6478 7642
rect 6502 7590 6516 7642
rect 6516 7590 6528 7642
rect 6528 7590 6558 7642
rect 6582 7590 6592 7642
rect 6592 7590 6638 7642
rect 6342 7588 6398 7590
rect 6422 7588 6478 7590
rect 6502 7588 6558 7590
rect 6582 7588 6638 7590
rect 5682 7098 5738 7100
rect 5762 7098 5818 7100
rect 5842 7098 5898 7100
rect 5922 7098 5978 7100
rect 5682 7046 5728 7098
rect 5728 7046 5738 7098
rect 5762 7046 5792 7098
rect 5792 7046 5804 7098
rect 5804 7046 5818 7098
rect 5842 7046 5856 7098
rect 5856 7046 5868 7098
rect 5868 7046 5898 7098
rect 5922 7046 5932 7098
rect 5932 7046 5978 7098
rect 5682 7044 5738 7046
rect 5762 7044 5818 7046
rect 5842 7044 5898 7046
rect 5922 7044 5978 7046
rect 5682 6010 5738 6012
rect 5762 6010 5818 6012
rect 5842 6010 5898 6012
rect 5922 6010 5978 6012
rect 5682 5958 5728 6010
rect 5728 5958 5738 6010
rect 5762 5958 5792 6010
rect 5792 5958 5804 6010
rect 5804 5958 5818 6010
rect 5842 5958 5856 6010
rect 5856 5958 5868 6010
rect 5868 5958 5898 6010
rect 5922 5958 5932 6010
rect 5932 5958 5978 6010
rect 5682 5956 5738 5958
rect 5762 5956 5818 5958
rect 5842 5956 5898 5958
rect 5922 5956 5978 5958
rect 3191 5466 3247 5468
rect 3271 5466 3327 5468
rect 3351 5466 3407 5468
rect 3431 5466 3487 5468
rect 3191 5414 3237 5466
rect 3237 5414 3247 5466
rect 3271 5414 3301 5466
rect 3301 5414 3313 5466
rect 3313 5414 3327 5466
rect 3351 5414 3365 5466
rect 3365 5414 3377 5466
rect 3377 5414 3407 5466
rect 3431 5414 3441 5466
rect 3441 5414 3487 5466
rect 3191 5412 3247 5414
rect 3271 5412 3327 5414
rect 3351 5412 3407 5414
rect 3431 5412 3487 5414
rect 2531 4922 2587 4924
rect 2611 4922 2667 4924
rect 2691 4922 2747 4924
rect 2771 4922 2827 4924
rect 2531 4870 2577 4922
rect 2577 4870 2587 4922
rect 2611 4870 2641 4922
rect 2641 4870 2653 4922
rect 2653 4870 2667 4922
rect 2691 4870 2705 4922
rect 2705 4870 2717 4922
rect 2717 4870 2747 4922
rect 2771 4870 2781 4922
rect 2781 4870 2827 4922
rect 2531 4868 2587 4870
rect 2611 4868 2667 4870
rect 2691 4868 2747 4870
rect 2771 4868 2827 4870
rect 3191 4378 3247 4380
rect 3271 4378 3327 4380
rect 3351 4378 3407 4380
rect 3431 4378 3487 4380
rect 3191 4326 3237 4378
rect 3237 4326 3247 4378
rect 3271 4326 3301 4378
rect 3301 4326 3313 4378
rect 3313 4326 3327 4378
rect 3351 4326 3365 4378
rect 3365 4326 3377 4378
rect 3377 4326 3407 4378
rect 3431 4326 3441 4378
rect 3441 4326 3487 4378
rect 3191 4324 3247 4326
rect 3271 4324 3327 4326
rect 3351 4324 3407 4326
rect 3431 4324 3487 4326
rect 2531 3834 2587 3836
rect 2611 3834 2667 3836
rect 2691 3834 2747 3836
rect 2771 3834 2827 3836
rect 2531 3782 2577 3834
rect 2577 3782 2587 3834
rect 2611 3782 2641 3834
rect 2641 3782 2653 3834
rect 2653 3782 2667 3834
rect 2691 3782 2705 3834
rect 2705 3782 2717 3834
rect 2717 3782 2747 3834
rect 2771 3782 2781 3834
rect 2781 3782 2827 3834
rect 2531 3780 2587 3782
rect 2611 3780 2667 3782
rect 2691 3780 2747 3782
rect 2771 3780 2827 3782
rect 846 3612 848 3632
rect 848 3612 900 3632
rect 900 3612 902 3632
rect 846 3576 902 3612
rect 3191 3290 3247 3292
rect 3271 3290 3327 3292
rect 3351 3290 3407 3292
rect 3431 3290 3487 3292
rect 3191 3238 3237 3290
rect 3237 3238 3247 3290
rect 3271 3238 3301 3290
rect 3301 3238 3313 3290
rect 3313 3238 3327 3290
rect 3351 3238 3365 3290
rect 3365 3238 3377 3290
rect 3377 3238 3407 3290
rect 3431 3238 3441 3290
rect 3441 3238 3487 3290
rect 3191 3236 3247 3238
rect 3271 3236 3327 3238
rect 3351 3236 3407 3238
rect 3431 3236 3487 3238
rect 846 2932 848 2952
rect 848 2932 900 2952
rect 900 2932 902 2952
rect 846 2896 902 2932
rect 2531 2746 2587 2748
rect 2611 2746 2667 2748
rect 2691 2746 2747 2748
rect 2771 2746 2827 2748
rect 2531 2694 2577 2746
rect 2577 2694 2587 2746
rect 2611 2694 2641 2746
rect 2641 2694 2653 2746
rect 2653 2694 2667 2746
rect 2691 2694 2705 2746
rect 2705 2694 2717 2746
rect 2717 2694 2747 2746
rect 2771 2694 2781 2746
rect 2781 2694 2827 2746
rect 2531 2692 2587 2694
rect 2611 2692 2667 2694
rect 2691 2692 2747 2694
rect 2771 2692 2827 2694
rect 6342 6554 6398 6556
rect 6422 6554 6478 6556
rect 6502 6554 6558 6556
rect 6582 6554 6638 6556
rect 6342 6502 6388 6554
rect 6388 6502 6398 6554
rect 6422 6502 6452 6554
rect 6452 6502 6464 6554
rect 6464 6502 6478 6554
rect 6502 6502 6516 6554
rect 6516 6502 6528 6554
rect 6528 6502 6558 6554
rect 6582 6502 6592 6554
rect 6592 6502 6638 6554
rect 6342 6500 6398 6502
rect 6422 6500 6478 6502
rect 6502 6500 6558 6502
rect 6582 6500 6638 6502
rect 9493 13082 9549 13084
rect 9573 13082 9629 13084
rect 9653 13082 9709 13084
rect 9733 13082 9789 13084
rect 9493 13030 9539 13082
rect 9539 13030 9549 13082
rect 9573 13030 9603 13082
rect 9603 13030 9615 13082
rect 9615 13030 9629 13082
rect 9653 13030 9667 13082
rect 9667 13030 9679 13082
rect 9679 13030 9709 13082
rect 9733 13030 9743 13082
rect 9743 13030 9789 13082
rect 9493 13028 9549 13030
rect 9573 13028 9629 13030
rect 9653 13028 9709 13030
rect 9733 13028 9789 13030
rect 8833 12538 8889 12540
rect 8913 12538 8969 12540
rect 8993 12538 9049 12540
rect 9073 12538 9129 12540
rect 8833 12486 8879 12538
rect 8879 12486 8889 12538
rect 8913 12486 8943 12538
rect 8943 12486 8955 12538
rect 8955 12486 8969 12538
rect 8993 12486 9007 12538
rect 9007 12486 9019 12538
rect 9019 12486 9049 12538
rect 9073 12486 9083 12538
rect 9083 12486 9129 12538
rect 8833 12484 8889 12486
rect 8913 12484 8969 12486
rect 8993 12484 9049 12486
rect 9073 12484 9129 12486
rect 7654 8472 7710 8528
rect 13358 13640 13414 13696
rect 11984 13626 12040 13628
rect 12064 13626 12120 13628
rect 12144 13626 12200 13628
rect 12224 13626 12280 13628
rect 11984 13574 12030 13626
rect 12030 13574 12040 13626
rect 12064 13574 12094 13626
rect 12094 13574 12106 13626
rect 12106 13574 12120 13626
rect 12144 13574 12158 13626
rect 12158 13574 12170 13626
rect 12170 13574 12200 13626
rect 12224 13574 12234 13626
rect 12234 13574 12280 13626
rect 11984 13572 12040 13574
rect 12064 13572 12120 13574
rect 12144 13572 12200 13574
rect 12224 13572 12280 13574
rect 12644 13082 12700 13084
rect 12724 13082 12780 13084
rect 12804 13082 12860 13084
rect 12884 13082 12940 13084
rect 12644 13030 12690 13082
rect 12690 13030 12700 13082
rect 12724 13030 12754 13082
rect 12754 13030 12766 13082
rect 12766 13030 12780 13082
rect 12804 13030 12818 13082
rect 12818 13030 12830 13082
rect 12830 13030 12860 13082
rect 12884 13030 12894 13082
rect 12894 13030 12940 13082
rect 12644 13028 12700 13030
rect 12724 13028 12780 13030
rect 12804 13028 12860 13030
rect 12884 13028 12940 13030
rect 13358 12960 13414 13016
rect 8833 11450 8889 11452
rect 8913 11450 8969 11452
rect 8993 11450 9049 11452
rect 9073 11450 9129 11452
rect 8833 11398 8879 11450
rect 8879 11398 8889 11450
rect 8913 11398 8943 11450
rect 8943 11398 8955 11450
rect 8955 11398 8969 11450
rect 8993 11398 9007 11450
rect 9007 11398 9019 11450
rect 9019 11398 9049 11450
rect 9073 11398 9083 11450
rect 9083 11398 9129 11450
rect 8833 11396 8889 11398
rect 8913 11396 8969 11398
rect 8993 11396 9049 11398
rect 9073 11396 9129 11398
rect 9493 11994 9549 11996
rect 9573 11994 9629 11996
rect 9653 11994 9709 11996
rect 9733 11994 9789 11996
rect 9493 11942 9539 11994
rect 9539 11942 9549 11994
rect 9573 11942 9603 11994
rect 9603 11942 9615 11994
rect 9615 11942 9629 11994
rect 9653 11942 9667 11994
rect 9667 11942 9679 11994
rect 9679 11942 9709 11994
rect 9733 11942 9743 11994
rect 9743 11942 9789 11994
rect 9493 11940 9549 11942
rect 9573 11940 9629 11942
rect 9653 11940 9709 11942
rect 9733 11940 9789 11942
rect 9493 10906 9549 10908
rect 9573 10906 9629 10908
rect 9653 10906 9709 10908
rect 9733 10906 9789 10908
rect 9493 10854 9539 10906
rect 9539 10854 9549 10906
rect 9573 10854 9603 10906
rect 9603 10854 9615 10906
rect 9615 10854 9629 10906
rect 9653 10854 9667 10906
rect 9667 10854 9679 10906
rect 9679 10854 9709 10906
rect 9733 10854 9743 10906
rect 9743 10854 9789 10906
rect 9493 10852 9549 10854
rect 9573 10852 9629 10854
rect 9653 10852 9709 10854
rect 9733 10852 9789 10854
rect 8833 10362 8889 10364
rect 8913 10362 8969 10364
rect 8993 10362 9049 10364
rect 9073 10362 9129 10364
rect 8833 10310 8879 10362
rect 8879 10310 8889 10362
rect 8913 10310 8943 10362
rect 8943 10310 8955 10362
rect 8955 10310 8969 10362
rect 8993 10310 9007 10362
rect 9007 10310 9019 10362
rect 9019 10310 9049 10362
rect 9073 10310 9083 10362
rect 9083 10310 9129 10362
rect 8833 10308 8889 10310
rect 8913 10308 8969 10310
rect 8993 10308 9049 10310
rect 9073 10308 9129 10310
rect 6342 5466 6398 5468
rect 6422 5466 6478 5468
rect 6502 5466 6558 5468
rect 6582 5466 6638 5468
rect 6342 5414 6388 5466
rect 6388 5414 6398 5466
rect 6422 5414 6452 5466
rect 6452 5414 6464 5466
rect 6464 5414 6478 5466
rect 6502 5414 6516 5466
rect 6516 5414 6528 5466
rect 6528 5414 6558 5466
rect 6582 5414 6592 5466
rect 6592 5414 6638 5466
rect 6342 5412 6398 5414
rect 6422 5412 6478 5414
rect 6502 5412 6558 5414
rect 6582 5412 6638 5414
rect 5682 4922 5738 4924
rect 5762 4922 5818 4924
rect 5842 4922 5898 4924
rect 5922 4922 5978 4924
rect 5682 4870 5728 4922
rect 5728 4870 5738 4922
rect 5762 4870 5792 4922
rect 5792 4870 5804 4922
rect 5804 4870 5818 4922
rect 5842 4870 5856 4922
rect 5856 4870 5868 4922
rect 5868 4870 5898 4922
rect 5922 4870 5932 4922
rect 5932 4870 5978 4922
rect 5682 4868 5738 4870
rect 5762 4868 5818 4870
rect 5842 4868 5898 4870
rect 5922 4868 5978 4870
rect 5682 3834 5738 3836
rect 5762 3834 5818 3836
rect 5842 3834 5898 3836
rect 5922 3834 5978 3836
rect 5682 3782 5728 3834
rect 5728 3782 5738 3834
rect 5762 3782 5792 3834
rect 5792 3782 5804 3834
rect 5804 3782 5818 3834
rect 5842 3782 5856 3834
rect 5856 3782 5868 3834
rect 5868 3782 5898 3834
rect 5922 3782 5932 3834
rect 5932 3782 5978 3834
rect 5682 3780 5738 3782
rect 5762 3780 5818 3782
rect 5842 3780 5898 3782
rect 5922 3780 5978 3782
rect 6342 4378 6398 4380
rect 6422 4378 6478 4380
rect 6502 4378 6558 4380
rect 6582 4378 6638 4380
rect 6342 4326 6388 4378
rect 6388 4326 6398 4378
rect 6422 4326 6452 4378
rect 6452 4326 6464 4378
rect 6464 4326 6478 4378
rect 6502 4326 6516 4378
rect 6516 4326 6528 4378
rect 6528 4326 6558 4378
rect 6582 4326 6592 4378
rect 6592 4326 6638 4378
rect 6342 4324 6398 4326
rect 6422 4324 6478 4326
rect 6502 4324 6558 4326
rect 6582 4324 6638 4326
rect 6342 3290 6398 3292
rect 6422 3290 6478 3292
rect 6502 3290 6558 3292
rect 6582 3290 6638 3292
rect 6342 3238 6388 3290
rect 6388 3238 6398 3290
rect 6422 3238 6452 3290
rect 6452 3238 6464 3290
rect 6464 3238 6478 3290
rect 6502 3238 6516 3290
rect 6516 3238 6528 3290
rect 6528 3238 6558 3290
rect 6582 3238 6592 3290
rect 6592 3238 6638 3290
rect 6342 3236 6398 3238
rect 6422 3236 6478 3238
rect 6502 3236 6558 3238
rect 6582 3236 6638 3238
rect 5682 2746 5738 2748
rect 5762 2746 5818 2748
rect 5842 2746 5898 2748
rect 5922 2746 5978 2748
rect 5682 2694 5728 2746
rect 5728 2694 5738 2746
rect 5762 2694 5792 2746
rect 5792 2694 5804 2746
rect 5804 2694 5818 2746
rect 5842 2694 5856 2746
rect 5856 2694 5868 2746
rect 5868 2694 5898 2746
rect 5922 2694 5932 2746
rect 5932 2694 5978 2746
rect 5682 2692 5738 2694
rect 5762 2692 5818 2694
rect 5842 2692 5898 2694
rect 5922 2692 5978 2694
rect 8833 9274 8889 9276
rect 8913 9274 8969 9276
rect 8993 9274 9049 9276
rect 9073 9274 9129 9276
rect 8833 9222 8879 9274
rect 8879 9222 8889 9274
rect 8913 9222 8943 9274
rect 8943 9222 8955 9274
rect 8955 9222 8969 9274
rect 8993 9222 9007 9274
rect 9007 9222 9019 9274
rect 9019 9222 9049 9274
rect 9073 9222 9083 9274
rect 9083 9222 9129 9274
rect 8833 9220 8889 9222
rect 8913 9220 8969 9222
rect 8993 9220 9049 9222
rect 9073 9220 9129 9222
rect 9493 9818 9549 9820
rect 9573 9818 9629 9820
rect 9653 9818 9709 9820
rect 9733 9818 9789 9820
rect 9493 9766 9539 9818
rect 9539 9766 9549 9818
rect 9573 9766 9603 9818
rect 9603 9766 9615 9818
rect 9615 9766 9629 9818
rect 9653 9766 9667 9818
rect 9667 9766 9679 9818
rect 9679 9766 9709 9818
rect 9733 9766 9743 9818
rect 9743 9766 9789 9818
rect 9493 9764 9549 9766
rect 9573 9764 9629 9766
rect 9653 9764 9709 9766
rect 9733 9764 9789 9766
rect 11984 12538 12040 12540
rect 12064 12538 12120 12540
rect 12144 12538 12200 12540
rect 12224 12538 12280 12540
rect 11984 12486 12030 12538
rect 12030 12486 12040 12538
rect 12064 12486 12094 12538
rect 12094 12486 12106 12538
rect 12106 12486 12120 12538
rect 12144 12486 12158 12538
rect 12158 12486 12170 12538
rect 12170 12486 12200 12538
rect 12224 12486 12234 12538
rect 12234 12486 12280 12538
rect 11984 12484 12040 12486
rect 12064 12484 12120 12486
rect 12144 12484 12200 12486
rect 12224 12484 12280 12486
rect 12644 11994 12700 11996
rect 12724 11994 12780 11996
rect 12804 11994 12860 11996
rect 12884 11994 12940 11996
rect 12644 11942 12690 11994
rect 12690 11942 12700 11994
rect 12724 11942 12754 11994
rect 12754 11942 12766 11994
rect 12766 11942 12780 11994
rect 12804 11942 12818 11994
rect 12818 11942 12830 11994
rect 12830 11942 12860 11994
rect 12884 11942 12894 11994
rect 12894 11942 12940 11994
rect 12644 11940 12700 11942
rect 12724 11940 12780 11942
rect 12804 11940 12860 11942
rect 12884 11940 12940 11942
rect 11984 11450 12040 11452
rect 12064 11450 12120 11452
rect 12144 11450 12200 11452
rect 12224 11450 12280 11452
rect 11984 11398 12030 11450
rect 12030 11398 12040 11450
rect 12064 11398 12094 11450
rect 12094 11398 12106 11450
rect 12106 11398 12120 11450
rect 12144 11398 12158 11450
rect 12158 11398 12170 11450
rect 12170 11398 12200 11450
rect 12224 11398 12234 11450
rect 12234 11398 12280 11450
rect 11984 11396 12040 11398
rect 12064 11396 12120 11398
rect 12144 11396 12200 11398
rect 12224 11396 12280 11398
rect 9493 8730 9549 8732
rect 9573 8730 9629 8732
rect 9653 8730 9709 8732
rect 9733 8730 9789 8732
rect 9493 8678 9539 8730
rect 9539 8678 9549 8730
rect 9573 8678 9603 8730
rect 9603 8678 9615 8730
rect 9615 8678 9629 8730
rect 9653 8678 9667 8730
rect 9667 8678 9679 8730
rect 9679 8678 9709 8730
rect 9733 8678 9743 8730
rect 9743 8678 9789 8730
rect 9493 8676 9549 8678
rect 9573 8676 9629 8678
rect 9653 8676 9709 8678
rect 9733 8676 9789 8678
rect 8666 8492 8722 8528
rect 8666 8472 8668 8492
rect 8668 8472 8720 8492
rect 8720 8472 8722 8492
rect 8833 8186 8889 8188
rect 8913 8186 8969 8188
rect 8993 8186 9049 8188
rect 9073 8186 9129 8188
rect 8833 8134 8879 8186
rect 8879 8134 8889 8186
rect 8913 8134 8943 8186
rect 8943 8134 8955 8186
rect 8955 8134 8969 8186
rect 8993 8134 9007 8186
rect 9007 8134 9019 8186
rect 9019 8134 9049 8186
rect 9073 8134 9083 8186
rect 9083 8134 9129 8186
rect 8833 8132 8889 8134
rect 8913 8132 8969 8134
rect 8993 8132 9049 8134
rect 9073 8132 9129 8134
rect 9493 7642 9549 7644
rect 9573 7642 9629 7644
rect 9653 7642 9709 7644
rect 9733 7642 9789 7644
rect 9493 7590 9539 7642
rect 9539 7590 9549 7642
rect 9573 7590 9603 7642
rect 9603 7590 9615 7642
rect 9615 7590 9629 7642
rect 9653 7590 9667 7642
rect 9667 7590 9679 7642
rect 9679 7590 9709 7642
rect 9733 7590 9743 7642
rect 9743 7590 9789 7642
rect 9493 7588 9549 7590
rect 9573 7588 9629 7590
rect 9653 7588 9709 7590
rect 9733 7588 9789 7590
rect 8574 6296 8630 6352
rect 8833 7098 8889 7100
rect 8913 7098 8969 7100
rect 8993 7098 9049 7100
rect 9073 7098 9129 7100
rect 8833 7046 8879 7098
rect 8879 7046 8889 7098
rect 8913 7046 8943 7098
rect 8943 7046 8955 7098
rect 8955 7046 8969 7098
rect 8993 7046 9007 7098
rect 9007 7046 9019 7098
rect 9019 7046 9049 7098
rect 9073 7046 9083 7098
rect 9083 7046 9129 7098
rect 8833 7044 8889 7046
rect 8913 7044 8969 7046
rect 8993 7044 9049 7046
rect 9073 7044 9129 7046
rect 9493 6554 9549 6556
rect 9573 6554 9629 6556
rect 9653 6554 9709 6556
rect 9733 6554 9789 6556
rect 9493 6502 9539 6554
rect 9539 6502 9549 6554
rect 9573 6502 9603 6554
rect 9603 6502 9615 6554
rect 9615 6502 9629 6554
rect 9653 6502 9667 6554
rect 9667 6502 9679 6554
rect 9679 6502 9709 6554
rect 9733 6502 9743 6554
rect 9743 6502 9789 6554
rect 9493 6500 9549 6502
rect 9573 6500 9629 6502
rect 9653 6500 9709 6502
rect 9733 6500 9789 6502
rect 9586 6316 9642 6352
rect 9586 6296 9588 6316
rect 9588 6296 9640 6316
rect 9640 6296 9642 6316
rect 8850 6160 8906 6216
rect 8833 6010 8889 6012
rect 8913 6010 8969 6012
rect 8993 6010 9049 6012
rect 9073 6010 9129 6012
rect 8833 5958 8879 6010
rect 8879 5958 8889 6010
rect 8913 5958 8943 6010
rect 8943 5958 8955 6010
rect 8955 5958 8969 6010
rect 8993 5958 9007 6010
rect 9007 5958 9019 6010
rect 9019 5958 9049 6010
rect 9073 5958 9083 6010
rect 9083 5958 9129 6010
rect 8833 5956 8889 5958
rect 8913 5956 8969 5958
rect 8993 5956 9049 5958
rect 9073 5956 9129 5958
rect 8833 4922 8889 4924
rect 8913 4922 8969 4924
rect 8993 4922 9049 4924
rect 9073 4922 9129 4924
rect 8833 4870 8879 4922
rect 8879 4870 8889 4922
rect 8913 4870 8943 4922
rect 8943 4870 8955 4922
rect 8955 4870 8969 4922
rect 8993 4870 9007 4922
rect 9007 4870 9019 4922
rect 9019 4870 9049 4922
rect 9073 4870 9083 4922
rect 9083 4870 9129 4922
rect 8833 4868 8889 4870
rect 8913 4868 8969 4870
rect 8993 4868 9049 4870
rect 9073 4868 9129 4870
rect 10230 6160 10286 6216
rect 12644 10906 12700 10908
rect 12724 10906 12780 10908
rect 12804 10906 12860 10908
rect 12884 10906 12940 10908
rect 12644 10854 12690 10906
rect 12690 10854 12700 10906
rect 12724 10854 12754 10906
rect 12754 10854 12766 10906
rect 12766 10854 12780 10906
rect 12804 10854 12818 10906
rect 12818 10854 12830 10906
rect 12830 10854 12860 10906
rect 12884 10854 12894 10906
rect 12894 10854 12940 10906
rect 12644 10852 12700 10854
rect 12724 10852 12780 10854
rect 12804 10852 12860 10854
rect 12884 10852 12940 10854
rect 11984 10362 12040 10364
rect 12064 10362 12120 10364
rect 12144 10362 12200 10364
rect 12224 10362 12280 10364
rect 11984 10310 12030 10362
rect 12030 10310 12040 10362
rect 12064 10310 12094 10362
rect 12094 10310 12106 10362
rect 12106 10310 12120 10362
rect 12144 10310 12158 10362
rect 12158 10310 12170 10362
rect 12170 10310 12200 10362
rect 12224 10310 12234 10362
rect 12234 10310 12280 10362
rect 11984 10308 12040 10310
rect 12064 10308 12120 10310
rect 12144 10308 12200 10310
rect 12224 10308 12280 10310
rect 12644 9818 12700 9820
rect 12724 9818 12780 9820
rect 12804 9818 12860 9820
rect 12884 9818 12940 9820
rect 12644 9766 12690 9818
rect 12690 9766 12700 9818
rect 12724 9766 12754 9818
rect 12754 9766 12766 9818
rect 12766 9766 12780 9818
rect 12804 9766 12818 9818
rect 12818 9766 12830 9818
rect 12830 9766 12860 9818
rect 12884 9766 12894 9818
rect 12894 9766 12940 9818
rect 12644 9764 12700 9766
rect 12724 9764 12780 9766
rect 12804 9764 12860 9766
rect 12884 9764 12940 9766
rect 11984 9274 12040 9276
rect 12064 9274 12120 9276
rect 12144 9274 12200 9276
rect 12224 9274 12280 9276
rect 11984 9222 12030 9274
rect 12030 9222 12040 9274
rect 12064 9222 12094 9274
rect 12094 9222 12106 9274
rect 12106 9222 12120 9274
rect 12144 9222 12158 9274
rect 12158 9222 12170 9274
rect 12170 9222 12200 9274
rect 12224 9222 12234 9274
rect 12234 9222 12280 9274
rect 11984 9220 12040 9222
rect 12064 9220 12120 9222
rect 12144 9220 12200 9222
rect 12224 9220 12280 9222
rect 11984 8186 12040 8188
rect 12064 8186 12120 8188
rect 12144 8186 12200 8188
rect 12224 8186 12280 8188
rect 11984 8134 12030 8186
rect 12030 8134 12040 8186
rect 12064 8134 12094 8186
rect 12094 8134 12106 8186
rect 12106 8134 12120 8186
rect 12144 8134 12158 8186
rect 12158 8134 12170 8186
rect 12170 8134 12200 8186
rect 12224 8134 12234 8186
rect 12234 8134 12280 8186
rect 11984 8132 12040 8134
rect 12064 8132 12120 8134
rect 12144 8132 12200 8134
rect 12224 8132 12280 8134
rect 12644 8730 12700 8732
rect 12724 8730 12780 8732
rect 12804 8730 12860 8732
rect 12884 8730 12940 8732
rect 12644 8678 12690 8730
rect 12690 8678 12700 8730
rect 12724 8678 12754 8730
rect 12754 8678 12766 8730
rect 12766 8678 12780 8730
rect 12804 8678 12818 8730
rect 12818 8678 12830 8730
rect 12830 8678 12860 8730
rect 12884 8678 12894 8730
rect 12894 8678 12940 8730
rect 12644 8676 12700 8678
rect 12724 8676 12780 8678
rect 12804 8676 12860 8678
rect 12884 8676 12940 8678
rect 12644 7642 12700 7644
rect 12724 7642 12780 7644
rect 12804 7642 12860 7644
rect 12884 7642 12940 7644
rect 12644 7590 12690 7642
rect 12690 7590 12700 7642
rect 12724 7590 12754 7642
rect 12754 7590 12766 7642
rect 12766 7590 12780 7642
rect 12804 7590 12818 7642
rect 12818 7590 12830 7642
rect 12830 7590 12860 7642
rect 12884 7590 12894 7642
rect 12894 7590 12940 7642
rect 12644 7588 12700 7590
rect 12724 7588 12780 7590
rect 12804 7588 12860 7590
rect 12884 7588 12940 7590
rect 11984 7098 12040 7100
rect 12064 7098 12120 7100
rect 12144 7098 12200 7100
rect 12224 7098 12280 7100
rect 11984 7046 12030 7098
rect 12030 7046 12040 7098
rect 12064 7046 12094 7098
rect 12094 7046 12106 7098
rect 12106 7046 12120 7098
rect 12144 7046 12158 7098
rect 12158 7046 12170 7098
rect 12170 7046 12200 7098
rect 12224 7046 12234 7098
rect 12234 7046 12280 7098
rect 11984 7044 12040 7046
rect 12064 7044 12120 7046
rect 12144 7044 12200 7046
rect 12224 7044 12280 7046
rect 12644 6554 12700 6556
rect 12724 6554 12780 6556
rect 12804 6554 12860 6556
rect 12884 6554 12940 6556
rect 12644 6502 12690 6554
rect 12690 6502 12700 6554
rect 12724 6502 12754 6554
rect 12754 6502 12766 6554
rect 12766 6502 12780 6554
rect 12804 6502 12818 6554
rect 12818 6502 12830 6554
rect 12830 6502 12860 6554
rect 12884 6502 12894 6554
rect 12894 6502 12940 6554
rect 12644 6500 12700 6502
rect 12724 6500 12780 6502
rect 12804 6500 12860 6502
rect 12884 6500 12940 6502
rect 9493 5466 9549 5468
rect 9573 5466 9629 5468
rect 9653 5466 9709 5468
rect 9733 5466 9789 5468
rect 9493 5414 9539 5466
rect 9539 5414 9549 5466
rect 9573 5414 9603 5466
rect 9603 5414 9615 5466
rect 9615 5414 9629 5466
rect 9653 5414 9667 5466
rect 9667 5414 9679 5466
rect 9679 5414 9709 5466
rect 9733 5414 9743 5466
rect 9743 5414 9789 5466
rect 9493 5412 9549 5414
rect 9573 5412 9629 5414
rect 9653 5412 9709 5414
rect 9733 5412 9789 5414
rect 11984 6010 12040 6012
rect 12064 6010 12120 6012
rect 12144 6010 12200 6012
rect 12224 6010 12280 6012
rect 11984 5958 12030 6010
rect 12030 5958 12040 6010
rect 12064 5958 12094 6010
rect 12094 5958 12106 6010
rect 12106 5958 12120 6010
rect 12144 5958 12158 6010
rect 12158 5958 12170 6010
rect 12170 5958 12200 6010
rect 12224 5958 12234 6010
rect 12234 5958 12280 6010
rect 11984 5956 12040 5958
rect 12064 5956 12120 5958
rect 12144 5956 12200 5958
rect 12224 5956 12280 5958
rect 12644 5466 12700 5468
rect 12724 5466 12780 5468
rect 12804 5466 12860 5468
rect 12884 5466 12940 5468
rect 12644 5414 12690 5466
rect 12690 5414 12700 5466
rect 12724 5414 12754 5466
rect 12754 5414 12766 5466
rect 12766 5414 12780 5466
rect 12804 5414 12818 5466
rect 12818 5414 12830 5466
rect 12830 5414 12860 5466
rect 12884 5414 12894 5466
rect 12894 5414 12940 5466
rect 12644 5412 12700 5414
rect 12724 5412 12780 5414
rect 12804 5412 12860 5414
rect 12884 5412 12940 5414
rect 8833 3834 8889 3836
rect 8913 3834 8969 3836
rect 8993 3834 9049 3836
rect 9073 3834 9129 3836
rect 8833 3782 8879 3834
rect 8879 3782 8889 3834
rect 8913 3782 8943 3834
rect 8943 3782 8955 3834
rect 8955 3782 8969 3834
rect 8993 3782 9007 3834
rect 9007 3782 9019 3834
rect 9019 3782 9049 3834
rect 9073 3782 9083 3834
rect 9083 3782 9129 3834
rect 8833 3780 8889 3782
rect 8913 3780 8969 3782
rect 8993 3780 9049 3782
rect 9073 3780 9129 3782
rect 9493 4378 9549 4380
rect 9573 4378 9629 4380
rect 9653 4378 9709 4380
rect 9733 4378 9789 4380
rect 9493 4326 9539 4378
rect 9539 4326 9549 4378
rect 9573 4326 9603 4378
rect 9603 4326 9615 4378
rect 9615 4326 9629 4378
rect 9653 4326 9667 4378
rect 9667 4326 9679 4378
rect 9679 4326 9709 4378
rect 9733 4326 9743 4378
rect 9743 4326 9789 4378
rect 9493 4324 9549 4326
rect 9573 4324 9629 4326
rect 9653 4324 9709 4326
rect 9733 4324 9789 4326
rect 9493 3290 9549 3292
rect 9573 3290 9629 3292
rect 9653 3290 9709 3292
rect 9733 3290 9789 3292
rect 9493 3238 9539 3290
rect 9539 3238 9549 3290
rect 9573 3238 9603 3290
rect 9603 3238 9615 3290
rect 9615 3238 9629 3290
rect 9653 3238 9667 3290
rect 9667 3238 9679 3290
rect 9679 3238 9709 3290
rect 9733 3238 9743 3290
rect 9743 3238 9789 3290
rect 9493 3236 9549 3238
rect 9573 3236 9629 3238
rect 9653 3236 9709 3238
rect 9733 3236 9789 3238
rect 11984 4922 12040 4924
rect 12064 4922 12120 4924
rect 12144 4922 12200 4924
rect 12224 4922 12280 4924
rect 11984 4870 12030 4922
rect 12030 4870 12040 4922
rect 12064 4870 12094 4922
rect 12094 4870 12106 4922
rect 12106 4870 12120 4922
rect 12144 4870 12158 4922
rect 12158 4870 12170 4922
rect 12170 4870 12200 4922
rect 12224 4870 12234 4922
rect 12234 4870 12280 4922
rect 11984 4868 12040 4870
rect 12064 4868 12120 4870
rect 12144 4868 12200 4870
rect 12224 4868 12280 4870
rect 8833 2746 8889 2748
rect 8913 2746 8969 2748
rect 8993 2746 9049 2748
rect 9073 2746 9129 2748
rect 8833 2694 8879 2746
rect 8879 2694 8889 2746
rect 8913 2694 8943 2746
rect 8943 2694 8955 2746
rect 8955 2694 8969 2746
rect 8993 2694 9007 2746
rect 9007 2694 9019 2746
rect 9019 2694 9049 2746
rect 9073 2694 9083 2746
rect 9083 2694 9129 2746
rect 8833 2692 8889 2694
rect 8913 2692 8969 2694
rect 8993 2692 9049 2694
rect 9073 2692 9129 2694
rect 11984 3834 12040 3836
rect 12064 3834 12120 3836
rect 12144 3834 12200 3836
rect 12224 3834 12280 3836
rect 11984 3782 12030 3834
rect 12030 3782 12040 3834
rect 12064 3782 12094 3834
rect 12094 3782 12106 3834
rect 12106 3782 12120 3834
rect 12144 3782 12158 3834
rect 12158 3782 12170 3834
rect 12170 3782 12200 3834
rect 12224 3782 12234 3834
rect 12234 3782 12280 3834
rect 11984 3780 12040 3782
rect 12064 3780 12120 3782
rect 12144 3780 12200 3782
rect 12224 3780 12280 3782
rect 12644 4378 12700 4380
rect 12724 4378 12780 4380
rect 12804 4378 12860 4380
rect 12884 4378 12940 4380
rect 12644 4326 12690 4378
rect 12690 4326 12700 4378
rect 12724 4326 12754 4378
rect 12754 4326 12766 4378
rect 12766 4326 12780 4378
rect 12804 4326 12818 4378
rect 12818 4326 12830 4378
rect 12830 4326 12860 4378
rect 12884 4326 12894 4378
rect 12894 4326 12940 4378
rect 12644 4324 12700 4326
rect 12724 4324 12780 4326
rect 12804 4324 12860 4326
rect 12884 4324 12940 4326
rect 13266 4120 13322 4176
rect 13358 3476 13360 3496
rect 13360 3476 13412 3496
rect 13412 3476 13414 3496
rect 13358 3440 13414 3476
rect 12644 3290 12700 3292
rect 12724 3290 12780 3292
rect 12804 3290 12860 3292
rect 12884 3290 12940 3292
rect 12644 3238 12690 3290
rect 12690 3238 12700 3290
rect 12724 3238 12754 3290
rect 12754 3238 12766 3290
rect 12766 3238 12780 3290
rect 12804 3238 12818 3290
rect 12818 3238 12830 3290
rect 12830 3238 12860 3290
rect 12884 3238 12894 3290
rect 12894 3238 12940 3290
rect 12644 3236 12700 3238
rect 12724 3236 12780 3238
rect 12804 3236 12860 3238
rect 12884 3236 12940 3238
rect 13358 2760 13414 2816
rect 11984 2746 12040 2748
rect 12064 2746 12120 2748
rect 12144 2746 12200 2748
rect 12224 2746 12280 2748
rect 11984 2694 12030 2746
rect 12030 2694 12040 2746
rect 12064 2694 12094 2746
rect 12094 2694 12106 2746
rect 12106 2694 12120 2746
rect 12144 2694 12158 2746
rect 12158 2694 12170 2746
rect 12170 2694 12200 2746
rect 12224 2694 12234 2746
rect 12234 2694 12280 2746
rect 11984 2692 12040 2694
rect 12064 2692 12120 2694
rect 12144 2692 12200 2694
rect 12224 2692 12280 2694
rect 3191 2202 3247 2204
rect 3271 2202 3327 2204
rect 3351 2202 3407 2204
rect 3431 2202 3487 2204
rect 3191 2150 3237 2202
rect 3237 2150 3247 2202
rect 3271 2150 3301 2202
rect 3301 2150 3313 2202
rect 3313 2150 3327 2202
rect 3351 2150 3365 2202
rect 3365 2150 3377 2202
rect 3377 2150 3407 2202
rect 3431 2150 3441 2202
rect 3441 2150 3487 2202
rect 3191 2148 3247 2150
rect 3271 2148 3327 2150
rect 3351 2148 3407 2150
rect 3431 2148 3487 2150
rect 6342 2202 6398 2204
rect 6422 2202 6478 2204
rect 6502 2202 6558 2204
rect 6582 2202 6638 2204
rect 6342 2150 6388 2202
rect 6388 2150 6398 2202
rect 6422 2150 6452 2202
rect 6452 2150 6464 2202
rect 6464 2150 6478 2202
rect 6502 2150 6516 2202
rect 6516 2150 6528 2202
rect 6528 2150 6558 2202
rect 6582 2150 6592 2202
rect 6592 2150 6638 2202
rect 6342 2148 6398 2150
rect 6422 2148 6478 2150
rect 6502 2148 6558 2150
rect 6582 2148 6638 2150
rect 9493 2202 9549 2204
rect 9573 2202 9629 2204
rect 9653 2202 9709 2204
rect 9733 2202 9789 2204
rect 9493 2150 9539 2202
rect 9539 2150 9549 2202
rect 9573 2150 9603 2202
rect 9603 2150 9615 2202
rect 9615 2150 9629 2202
rect 9653 2150 9667 2202
rect 9667 2150 9679 2202
rect 9679 2150 9709 2202
rect 9733 2150 9743 2202
rect 9743 2150 9789 2202
rect 9493 2148 9549 2150
rect 9573 2148 9629 2150
rect 9653 2148 9709 2150
rect 9733 2148 9789 2150
rect 12644 2202 12700 2204
rect 12724 2202 12780 2204
rect 12804 2202 12860 2204
rect 12884 2202 12940 2204
rect 12644 2150 12690 2202
rect 12690 2150 12700 2202
rect 12724 2150 12754 2202
rect 12754 2150 12766 2202
rect 12766 2150 12780 2202
rect 12804 2150 12818 2202
rect 12818 2150 12830 2202
rect 12830 2150 12860 2202
rect 12884 2150 12894 2202
rect 12894 2150 12940 2202
rect 12644 2148 12700 2150
rect 12724 2148 12780 2150
rect 12804 2148 12860 2150
rect 12884 2148 12940 2150
<< metal3 >>
rect 2521 14720 2837 14721
rect 2521 14656 2527 14720
rect 2591 14656 2607 14720
rect 2671 14656 2687 14720
rect 2751 14656 2767 14720
rect 2831 14656 2837 14720
rect 2521 14655 2837 14656
rect 5672 14720 5988 14721
rect 5672 14656 5678 14720
rect 5742 14656 5758 14720
rect 5822 14656 5838 14720
rect 5902 14656 5918 14720
rect 5982 14656 5988 14720
rect 5672 14655 5988 14656
rect 8823 14720 9139 14721
rect 8823 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9069 14720
rect 9133 14656 9139 14720
rect 8823 14655 9139 14656
rect 11974 14720 12290 14721
rect 11974 14656 11980 14720
rect 12044 14656 12060 14720
rect 12124 14656 12140 14720
rect 12204 14656 12220 14720
rect 12284 14656 12290 14720
rect 11974 14655 12290 14656
rect 3181 14176 3497 14177
rect 3181 14112 3187 14176
rect 3251 14112 3267 14176
rect 3331 14112 3347 14176
rect 3411 14112 3427 14176
rect 3491 14112 3497 14176
rect 3181 14111 3497 14112
rect 6332 14176 6648 14177
rect 6332 14112 6338 14176
rect 6402 14112 6418 14176
rect 6482 14112 6498 14176
rect 6562 14112 6578 14176
rect 6642 14112 6648 14176
rect 6332 14111 6648 14112
rect 9483 14176 9799 14177
rect 9483 14112 9489 14176
rect 9553 14112 9569 14176
rect 9633 14112 9649 14176
rect 9713 14112 9729 14176
rect 9793 14112 9799 14176
rect 9483 14111 9799 14112
rect 12634 14176 12950 14177
rect 12634 14112 12640 14176
rect 12704 14112 12720 14176
rect 12784 14112 12800 14176
rect 12864 14112 12880 14176
rect 12944 14112 12950 14176
rect 12634 14111 12950 14112
rect 0 13698 800 13728
rect 1393 13698 1459 13701
rect 0 13696 1459 13698
rect 0 13640 1398 13696
rect 1454 13640 1459 13696
rect 0 13638 1459 13640
rect 0 13608 800 13638
rect 1393 13635 1459 13638
rect 13353 13698 13419 13701
rect 14087 13698 14887 13728
rect 13353 13696 14887 13698
rect 13353 13640 13358 13696
rect 13414 13640 14887 13696
rect 13353 13638 14887 13640
rect 13353 13635 13419 13638
rect 2521 13632 2837 13633
rect 2521 13568 2527 13632
rect 2591 13568 2607 13632
rect 2671 13568 2687 13632
rect 2751 13568 2767 13632
rect 2831 13568 2837 13632
rect 2521 13567 2837 13568
rect 5672 13632 5988 13633
rect 5672 13568 5678 13632
rect 5742 13568 5758 13632
rect 5822 13568 5838 13632
rect 5902 13568 5918 13632
rect 5982 13568 5988 13632
rect 5672 13567 5988 13568
rect 8823 13632 9139 13633
rect 8823 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9069 13632
rect 9133 13568 9139 13632
rect 8823 13567 9139 13568
rect 11974 13632 12290 13633
rect 11974 13568 11980 13632
rect 12044 13568 12060 13632
rect 12124 13568 12140 13632
rect 12204 13568 12220 13632
rect 12284 13568 12290 13632
rect 14087 13608 14887 13638
rect 11974 13567 12290 13568
rect 841 13154 907 13157
rect 798 13152 907 13154
rect 798 13096 846 13152
rect 902 13096 907 13152
rect 798 13091 907 13096
rect 798 13048 858 13091
rect 0 12958 858 13048
rect 3181 13088 3497 13089
rect 3181 13024 3187 13088
rect 3251 13024 3267 13088
rect 3331 13024 3347 13088
rect 3411 13024 3427 13088
rect 3491 13024 3497 13088
rect 3181 13023 3497 13024
rect 6332 13088 6648 13089
rect 6332 13024 6338 13088
rect 6402 13024 6418 13088
rect 6482 13024 6498 13088
rect 6562 13024 6578 13088
rect 6642 13024 6648 13088
rect 6332 13023 6648 13024
rect 9483 13088 9799 13089
rect 9483 13024 9489 13088
rect 9553 13024 9569 13088
rect 9633 13024 9649 13088
rect 9713 13024 9729 13088
rect 9793 13024 9799 13088
rect 9483 13023 9799 13024
rect 12634 13088 12950 13089
rect 12634 13024 12640 13088
rect 12704 13024 12720 13088
rect 12784 13024 12800 13088
rect 12864 13024 12880 13088
rect 12944 13024 12950 13088
rect 12634 13023 12950 13024
rect 13353 13018 13419 13021
rect 14087 13018 14887 13048
rect 13353 13016 14887 13018
rect 13353 12960 13358 13016
rect 13414 12960 14887 13016
rect 13353 12958 14887 12960
rect 0 12928 800 12958
rect 13353 12955 13419 12958
rect 14087 12928 14887 12958
rect 2521 12544 2837 12545
rect 2521 12480 2527 12544
rect 2591 12480 2607 12544
rect 2671 12480 2687 12544
rect 2751 12480 2767 12544
rect 2831 12480 2837 12544
rect 2521 12479 2837 12480
rect 5672 12544 5988 12545
rect 5672 12480 5678 12544
rect 5742 12480 5758 12544
rect 5822 12480 5838 12544
rect 5902 12480 5918 12544
rect 5982 12480 5988 12544
rect 5672 12479 5988 12480
rect 8823 12544 9139 12545
rect 8823 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9069 12544
rect 9133 12480 9139 12544
rect 8823 12479 9139 12480
rect 11974 12544 12290 12545
rect 11974 12480 11980 12544
rect 12044 12480 12060 12544
rect 12124 12480 12140 12544
rect 12204 12480 12220 12544
rect 12284 12480 12290 12544
rect 11974 12479 12290 12480
rect 0 12338 800 12368
rect 6126 12338 6132 12340
rect 0 12278 6132 12338
rect 0 12248 800 12278
rect 6126 12276 6132 12278
rect 6196 12276 6202 12340
rect 3181 12000 3497 12001
rect 3181 11936 3187 12000
rect 3251 11936 3267 12000
rect 3331 11936 3347 12000
rect 3411 11936 3427 12000
rect 3491 11936 3497 12000
rect 3181 11935 3497 11936
rect 6332 12000 6648 12001
rect 6332 11936 6338 12000
rect 6402 11936 6418 12000
rect 6482 11936 6498 12000
rect 6562 11936 6578 12000
rect 6642 11936 6648 12000
rect 6332 11935 6648 11936
rect 9483 12000 9799 12001
rect 9483 11936 9489 12000
rect 9553 11936 9569 12000
rect 9633 11936 9649 12000
rect 9713 11936 9729 12000
rect 9793 11936 9799 12000
rect 9483 11935 9799 11936
rect 12634 12000 12950 12001
rect 12634 11936 12640 12000
rect 12704 11936 12720 12000
rect 12784 11936 12800 12000
rect 12864 11936 12880 12000
rect 12944 11936 12950 12000
rect 12634 11935 12950 11936
rect 2521 11456 2837 11457
rect 2521 11392 2527 11456
rect 2591 11392 2607 11456
rect 2671 11392 2687 11456
rect 2751 11392 2767 11456
rect 2831 11392 2837 11456
rect 2521 11391 2837 11392
rect 5672 11456 5988 11457
rect 5672 11392 5678 11456
rect 5742 11392 5758 11456
rect 5822 11392 5838 11456
rect 5902 11392 5918 11456
rect 5982 11392 5988 11456
rect 5672 11391 5988 11392
rect 8823 11456 9139 11457
rect 8823 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9069 11456
rect 9133 11392 9139 11456
rect 8823 11391 9139 11392
rect 11974 11456 12290 11457
rect 11974 11392 11980 11456
rect 12044 11392 12060 11456
rect 12124 11392 12140 11456
rect 12204 11392 12220 11456
rect 12284 11392 12290 11456
rect 11974 11391 12290 11392
rect 3181 10912 3497 10913
rect 3181 10848 3187 10912
rect 3251 10848 3267 10912
rect 3331 10848 3347 10912
rect 3411 10848 3427 10912
rect 3491 10848 3497 10912
rect 3181 10847 3497 10848
rect 6332 10912 6648 10913
rect 6332 10848 6338 10912
rect 6402 10848 6418 10912
rect 6482 10848 6498 10912
rect 6562 10848 6578 10912
rect 6642 10848 6648 10912
rect 6332 10847 6648 10848
rect 9483 10912 9799 10913
rect 9483 10848 9489 10912
rect 9553 10848 9569 10912
rect 9633 10848 9649 10912
rect 9713 10848 9729 10912
rect 9793 10848 9799 10912
rect 9483 10847 9799 10848
rect 12634 10912 12950 10913
rect 12634 10848 12640 10912
rect 12704 10848 12720 10912
rect 12784 10848 12800 10912
rect 12864 10848 12880 10912
rect 12944 10848 12950 10912
rect 12634 10847 12950 10848
rect 2521 10368 2837 10369
rect 2521 10304 2527 10368
rect 2591 10304 2607 10368
rect 2671 10304 2687 10368
rect 2751 10304 2767 10368
rect 2831 10304 2837 10368
rect 2521 10303 2837 10304
rect 5672 10368 5988 10369
rect 5672 10304 5678 10368
rect 5742 10304 5758 10368
rect 5822 10304 5838 10368
rect 5902 10304 5918 10368
rect 5982 10304 5988 10368
rect 5672 10303 5988 10304
rect 8823 10368 9139 10369
rect 8823 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9069 10368
rect 9133 10304 9139 10368
rect 8823 10303 9139 10304
rect 11974 10368 12290 10369
rect 11974 10304 11980 10368
rect 12044 10304 12060 10368
rect 12124 10304 12140 10368
rect 12204 10304 12220 10368
rect 12284 10304 12290 10368
rect 11974 10303 12290 10304
rect 3181 9824 3497 9825
rect 3181 9760 3187 9824
rect 3251 9760 3267 9824
rect 3331 9760 3347 9824
rect 3411 9760 3427 9824
rect 3491 9760 3497 9824
rect 3181 9759 3497 9760
rect 6332 9824 6648 9825
rect 6332 9760 6338 9824
rect 6402 9760 6418 9824
rect 6482 9760 6498 9824
rect 6562 9760 6578 9824
rect 6642 9760 6648 9824
rect 6332 9759 6648 9760
rect 9483 9824 9799 9825
rect 9483 9760 9489 9824
rect 9553 9760 9569 9824
rect 9633 9760 9649 9824
rect 9713 9760 9729 9824
rect 9793 9760 9799 9824
rect 9483 9759 9799 9760
rect 12634 9824 12950 9825
rect 12634 9760 12640 9824
rect 12704 9760 12720 9824
rect 12784 9760 12800 9824
rect 12864 9760 12880 9824
rect 12944 9760 12950 9824
rect 12634 9759 12950 9760
rect 6126 9556 6132 9620
rect 6196 9618 6202 9620
rect 6545 9618 6611 9621
rect 6196 9616 6611 9618
rect 6196 9560 6550 9616
rect 6606 9560 6611 9616
rect 6196 9558 6611 9560
rect 6196 9556 6202 9558
rect 6545 9555 6611 9558
rect 2521 9280 2837 9281
rect 2521 9216 2527 9280
rect 2591 9216 2607 9280
rect 2671 9216 2687 9280
rect 2751 9216 2767 9280
rect 2831 9216 2837 9280
rect 2521 9215 2837 9216
rect 5672 9280 5988 9281
rect 5672 9216 5678 9280
rect 5742 9216 5758 9280
rect 5822 9216 5838 9280
rect 5902 9216 5918 9280
rect 5982 9216 5988 9280
rect 5672 9215 5988 9216
rect 8823 9280 9139 9281
rect 8823 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9069 9280
rect 9133 9216 9139 9280
rect 8823 9215 9139 9216
rect 11974 9280 12290 9281
rect 11974 9216 11980 9280
rect 12044 9216 12060 9280
rect 12124 9216 12140 9280
rect 12204 9216 12220 9280
rect 12284 9216 12290 9280
rect 11974 9215 12290 9216
rect 3181 8736 3497 8737
rect 3181 8672 3187 8736
rect 3251 8672 3267 8736
rect 3331 8672 3347 8736
rect 3411 8672 3427 8736
rect 3491 8672 3497 8736
rect 3181 8671 3497 8672
rect 6332 8736 6648 8737
rect 6332 8672 6338 8736
rect 6402 8672 6418 8736
rect 6482 8672 6498 8736
rect 6562 8672 6578 8736
rect 6642 8672 6648 8736
rect 6332 8671 6648 8672
rect 9483 8736 9799 8737
rect 9483 8672 9489 8736
rect 9553 8672 9569 8736
rect 9633 8672 9649 8736
rect 9713 8672 9729 8736
rect 9793 8672 9799 8736
rect 9483 8671 9799 8672
rect 12634 8736 12950 8737
rect 12634 8672 12640 8736
rect 12704 8672 12720 8736
rect 12784 8672 12800 8736
rect 12864 8672 12880 8736
rect 12944 8672 12950 8736
rect 12634 8671 12950 8672
rect 7649 8530 7715 8533
rect 8661 8530 8727 8533
rect 7649 8528 8727 8530
rect 7649 8472 7654 8528
rect 7710 8472 8666 8528
rect 8722 8472 8727 8528
rect 7649 8470 8727 8472
rect 7649 8467 7715 8470
rect 8661 8467 8727 8470
rect 2521 8192 2837 8193
rect 2521 8128 2527 8192
rect 2591 8128 2607 8192
rect 2671 8128 2687 8192
rect 2751 8128 2767 8192
rect 2831 8128 2837 8192
rect 2521 8127 2837 8128
rect 5672 8192 5988 8193
rect 5672 8128 5678 8192
rect 5742 8128 5758 8192
rect 5822 8128 5838 8192
rect 5902 8128 5918 8192
rect 5982 8128 5988 8192
rect 5672 8127 5988 8128
rect 8823 8192 9139 8193
rect 8823 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9069 8192
rect 9133 8128 9139 8192
rect 8823 8127 9139 8128
rect 11974 8192 12290 8193
rect 11974 8128 11980 8192
rect 12044 8128 12060 8192
rect 12124 8128 12140 8192
rect 12204 8128 12220 8192
rect 12284 8128 12290 8192
rect 11974 8127 12290 8128
rect 3181 7648 3497 7649
rect 3181 7584 3187 7648
rect 3251 7584 3267 7648
rect 3331 7584 3347 7648
rect 3411 7584 3427 7648
rect 3491 7584 3497 7648
rect 3181 7583 3497 7584
rect 6332 7648 6648 7649
rect 6332 7584 6338 7648
rect 6402 7584 6418 7648
rect 6482 7584 6498 7648
rect 6562 7584 6578 7648
rect 6642 7584 6648 7648
rect 6332 7583 6648 7584
rect 9483 7648 9799 7649
rect 9483 7584 9489 7648
rect 9553 7584 9569 7648
rect 9633 7584 9649 7648
rect 9713 7584 9729 7648
rect 9793 7584 9799 7648
rect 9483 7583 9799 7584
rect 12634 7648 12950 7649
rect 12634 7584 12640 7648
rect 12704 7584 12720 7648
rect 12784 7584 12800 7648
rect 12864 7584 12880 7648
rect 12944 7584 12950 7648
rect 12634 7583 12950 7584
rect 2521 7104 2837 7105
rect 2521 7040 2527 7104
rect 2591 7040 2607 7104
rect 2671 7040 2687 7104
rect 2751 7040 2767 7104
rect 2831 7040 2837 7104
rect 2521 7039 2837 7040
rect 5672 7104 5988 7105
rect 5672 7040 5678 7104
rect 5742 7040 5758 7104
rect 5822 7040 5838 7104
rect 5902 7040 5918 7104
rect 5982 7040 5988 7104
rect 5672 7039 5988 7040
rect 8823 7104 9139 7105
rect 8823 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9069 7104
rect 9133 7040 9139 7104
rect 8823 7039 9139 7040
rect 11974 7104 12290 7105
rect 11974 7040 11980 7104
rect 12044 7040 12060 7104
rect 12124 7040 12140 7104
rect 12204 7040 12220 7104
rect 12284 7040 12290 7104
rect 11974 7039 12290 7040
rect 3181 6560 3497 6561
rect 3181 6496 3187 6560
rect 3251 6496 3267 6560
rect 3331 6496 3347 6560
rect 3411 6496 3427 6560
rect 3491 6496 3497 6560
rect 3181 6495 3497 6496
rect 6332 6560 6648 6561
rect 6332 6496 6338 6560
rect 6402 6496 6418 6560
rect 6482 6496 6498 6560
rect 6562 6496 6578 6560
rect 6642 6496 6648 6560
rect 6332 6495 6648 6496
rect 9483 6560 9799 6561
rect 9483 6496 9489 6560
rect 9553 6496 9569 6560
rect 9633 6496 9649 6560
rect 9713 6496 9729 6560
rect 9793 6496 9799 6560
rect 9483 6495 9799 6496
rect 12634 6560 12950 6561
rect 12634 6496 12640 6560
rect 12704 6496 12720 6560
rect 12784 6496 12800 6560
rect 12864 6496 12880 6560
rect 12944 6496 12950 6560
rect 12634 6495 12950 6496
rect 8569 6354 8635 6357
rect 9581 6354 9647 6357
rect 8569 6352 9647 6354
rect 8569 6296 8574 6352
rect 8630 6296 9586 6352
rect 9642 6296 9647 6352
rect 8569 6294 9647 6296
rect 8569 6291 8635 6294
rect 9581 6291 9647 6294
rect 8845 6218 8911 6221
rect 10225 6218 10291 6221
rect 8845 6216 10291 6218
rect 8845 6160 8850 6216
rect 8906 6160 10230 6216
rect 10286 6160 10291 6216
rect 8845 6158 10291 6160
rect 8845 6155 8911 6158
rect 10225 6155 10291 6158
rect 2521 6016 2837 6017
rect 2521 5952 2527 6016
rect 2591 5952 2607 6016
rect 2671 5952 2687 6016
rect 2751 5952 2767 6016
rect 2831 5952 2837 6016
rect 2521 5951 2837 5952
rect 5672 6016 5988 6017
rect 5672 5952 5678 6016
rect 5742 5952 5758 6016
rect 5822 5952 5838 6016
rect 5902 5952 5918 6016
rect 5982 5952 5988 6016
rect 5672 5951 5988 5952
rect 8823 6016 9139 6017
rect 8823 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9069 6016
rect 9133 5952 9139 6016
rect 8823 5951 9139 5952
rect 11974 6016 12290 6017
rect 11974 5952 11980 6016
rect 12044 5952 12060 6016
rect 12124 5952 12140 6016
rect 12204 5952 12220 6016
rect 12284 5952 12290 6016
rect 11974 5951 12290 5952
rect 3181 5472 3497 5473
rect 3181 5408 3187 5472
rect 3251 5408 3267 5472
rect 3331 5408 3347 5472
rect 3411 5408 3427 5472
rect 3491 5408 3497 5472
rect 3181 5407 3497 5408
rect 6332 5472 6648 5473
rect 6332 5408 6338 5472
rect 6402 5408 6418 5472
rect 6482 5408 6498 5472
rect 6562 5408 6578 5472
rect 6642 5408 6648 5472
rect 6332 5407 6648 5408
rect 9483 5472 9799 5473
rect 9483 5408 9489 5472
rect 9553 5408 9569 5472
rect 9633 5408 9649 5472
rect 9713 5408 9729 5472
rect 9793 5408 9799 5472
rect 9483 5407 9799 5408
rect 12634 5472 12950 5473
rect 12634 5408 12640 5472
rect 12704 5408 12720 5472
rect 12784 5408 12800 5472
rect 12864 5408 12880 5472
rect 12944 5408 12950 5472
rect 12634 5407 12950 5408
rect 2521 4928 2837 4929
rect 2521 4864 2527 4928
rect 2591 4864 2607 4928
rect 2671 4864 2687 4928
rect 2751 4864 2767 4928
rect 2831 4864 2837 4928
rect 2521 4863 2837 4864
rect 5672 4928 5988 4929
rect 5672 4864 5678 4928
rect 5742 4864 5758 4928
rect 5822 4864 5838 4928
rect 5902 4864 5918 4928
rect 5982 4864 5988 4928
rect 5672 4863 5988 4864
rect 8823 4928 9139 4929
rect 8823 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9069 4928
rect 9133 4864 9139 4928
rect 8823 4863 9139 4864
rect 11974 4928 12290 4929
rect 11974 4864 11980 4928
rect 12044 4864 12060 4928
rect 12124 4864 12140 4928
rect 12204 4864 12220 4928
rect 12284 4864 12290 4928
rect 11974 4863 12290 4864
rect 3181 4384 3497 4385
rect 3181 4320 3187 4384
rect 3251 4320 3267 4384
rect 3331 4320 3347 4384
rect 3411 4320 3427 4384
rect 3491 4320 3497 4384
rect 3181 4319 3497 4320
rect 6332 4384 6648 4385
rect 6332 4320 6338 4384
rect 6402 4320 6418 4384
rect 6482 4320 6498 4384
rect 6562 4320 6578 4384
rect 6642 4320 6648 4384
rect 6332 4319 6648 4320
rect 9483 4384 9799 4385
rect 9483 4320 9489 4384
rect 9553 4320 9569 4384
rect 9633 4320 9649 4384
rect 9713 4320 9729 4384
rect 9793 4320 9799 4384
rect 9483 4319 9799 4320
rect 12634 4384 12950 4385
rect 12634 4320 12640 4384
rect 12704 4320 12720 4384
rect 12784 4320 12800 4384
rect 12864 4320 12880 4384
rect 12944 4320 12950 4384
rect 12634 4319 12950 4320
rect 13261 4178 13327 4181
rect 14087 4178 14887 4208
rect 13261 4176 14887 4178
rect 13261 4120 13266 4176
rect 13322 4120 14887 4176
rect 13261 4118 14887 4120
rect 13261 4115 13327 4118
rect 14087 4088 14887 4118
rect 2521 3840 2837 3841
rect 2521 3776 2527 3840
rect 2591 3776 2607 3840
rect 2671 3776 2687 3840
rect 2751 3776 2767 3840
rect 2831 3776 2837 3840
rect 2521 3775 2837 3776
rect 5672 3840 5988 3841
rect 5672 3776 5678 3840
rect 5742 3776 5758 3840
rect 5822 3776 5838 3840
rect 5902 3776 5918 3840
rect 5982 3776 5988 3840
rect 5672 3775 5988 3776
rect 8823 3840 9139 3841
rect 8823 3776 8829 3840
rect 8893 3776 8909 3840
rect 8973 3776 8989 3840
rect 9053 3776 9069 3840
rect 9133 3776 9139 3840
rect 8823 3775 9139 3776
rect 11974 3840 12290 3841
rect 11974 3776 11980 3840
rect 12044 3776 12060 3840
rect 12124 3776 12140 3840
rect 12204 3776 12220 3840
rect 12284 3776 12290 3840
rect 11974 3775 12290 3776
rect 841 3634 907 3637
rect 798 3632 907 3634
rect 798 3576 846 3632
rect 902 3576 907 3632
rect 798 3571 907 3576
rect 798 3528 858 3571
rect 0 3438 858 3528
rect 13353 3498 13419 3501
rect 14087 3498 14887 3528
rect 13353 3496 14887 3498
rect 13353 3440 13358 3496
rect 13414 3440 14887 3496
rect 13353 3438 14887 3440
rect 0 3408 800 3438
rect 13353 3435 13419 3438
rect 14087 3408 14887 3438
rect 3181 3296 3497 3297
rect 3181 3232 3187 3296
rect 3251 3232 3267 3296
rect 3331 3232 3347 3296
rect 3411 3232 3427 3296
rect 3491 3232 3497 3296
rect 3181 3231 3497 3232
rect 6332 3296 6648 3297
rect 6332 3232 6338 3296
rect 6402 3232 6418 3296
rect 6482 3232 6498 3296
rect 6562 3232 6578 3296
rect 6642 3232 6648 3296
rect 6332 3231 6648 3232
rect 9483 3296 9799 3297
rect 9483 3232 9489 3296
rect 9553 3232 9569 3296
rect 9633 3232 9649 3296
rect 9713 3232 9729 3296
rect 9793 3232 9799 3296
rect 9483 3231 9799 3232
rect 12634 3296 12950 3297
rect 12634 3232 12640 3296
rect 12704 3232 12720 3296
rect 12784 3232 12800 3296
rect 12864 3232 12880 3296
rect 12944 3232 12950 3296
rect 12634 3231 12950 3232
rect 841 2954 907 2957
rect 798 2952 907 2954
rect 798 2896 846 2952
rect 902 2896 907 2952
rect 798 2891 907 2896
rect 798 2848 858 2891
rect 0 2758 858 2848
rect 13353 2818 13419 2821
rect 14087 2818 14887 2848
rect 13353 2816 14887 2818
rect 13353 2760 13358 2816
rect 13414 2760 14887 2816
rect 13353 2758 14887 2760
rect 0 2728 800 2758
rect 13353 2755 13419 2758
rect 2521 2752 2837 2753
rect 2521 2688 2527 2752
rect 2591 2688 2607 2752
rect 2671 2688 2687 2752
rect 2751 2688 2767 2752
rect 2831 2688 2837 2752
rect 2521 2687 2837 2688
rect 5672 2752 5988 2753
rect 5672 2688 5678 2752
rect 5742 2688 5758 2752
rect 5822 2688 5838 2752
rect 5902 2688 5918 2752
rect 5982 2688 5988 2752
rect 5672 2687 5988 2688
rect 8823 2752 9139 2753
rect 8823 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9069 2752
rect 9133 2688 9139 2752
rect 8823 2687 9139 2688
rect 11974 2752 12290 2753
rect 11974 2688 11980 2752
rect 12044 2688 12060 2752
rect 12124 2688 12140 2752
rect 12204 2688 12220 2752
rect 12284 2688 12290 2752
rect 14087 2728 14887 2758
rect 11974 2687 12290 2688
rect 3181 2208 3497 2209
rect 3181 2144 3187 2208
rect 3251 2144 3267 2208
rect 3331 2144 3347 2208
rect 3411 2144 3427 2208
rect 3491 2144 3497 2208
rect 3181 2143 3497 2144
rect 6332 2208 6648 2209
rect 6332 2144 6338 2208
rect 6402 2144 6418 2208
rect 6482 2144 6498 2208
rect 6562 2144 6578 2208
rect 6642 2144 6648 2208
rect 6332 2143 6648 2144
rect 9483 2208 9799 2209
rect 9483 2144 9489 2208
rect 9553 2144 9569 2208
rect 9633 2144 9649 2208
rect 9713 2144 9729 2208
rect 9793 2144 9799 2208
rect 9483 2143 9799 2144
rect 12634 2208 12950 2209
rect 12634 2144 12640 2208
rect 12704 2144 12720 2208
rect 12784 2144 12800 2208
rect 12864 2144 12880 2208
rect 12944 2144 12950 2208
rect 12634 2143 12950 2144
<< via3 >>
rect 2527 14716 2591 14720
rect 2527 14660 2531 14716
rect 2531 14660 2587 14716
rect 2587 14660 2591 14716
rect 2527 14656 2591 14660
rect 2607 14716 2671 14720
rect 2607 14660 2611 14716
rect 2611 14660 2667 14716
rect 2667 14660 2671 14716
rect 2607 14656 2671 14660
rect 2687 14716 2751 14720
rect 2687 14660 2691 14716
rect 2691 14660 2747 14716
rect 2747 14660 2751 14716
rect 2687 14656 2751 14660
rect 2767 14716 2831 14720
rect 2767 14660 2771 14716
rect 2771 14660 2827 14716
rect 2827 14660 2831 14716
rect 2767 14656 2831 14660
rect 5678 14716 5742 14720
rect 5678 14660 5682 14716
rect 5682 14660 5738 14716
rect 5738 14660 5742 14716
rect 5678 14656 5742 14660
rect 5758 14716 5822 14720
rect 5758 14660 5762 14716
rect 5762 14660 5818 14716
rect 5818 14660 5822 14716
rect 5758 14656 5822 14660
rect 5838 14716 5902 14720
rect 5838 14660 5842 14716
rect 5842 14660 5898 14716
rect 5898 14660 5902 14716
rect 5838 14656 5902 14660
rect 5918 14716 5982 14720
rect 5918 14660 5922 14716
rect 5922 14660 5978 14716
rect 5978 14660 5982 14716
rect 5918 14656 5982 14660
rect 8829 14716 8893 14720
rect 8829 14660 8833 14716
rect 8833 14660 8889 14716
rect 8889 14660 8893 14716
rect 8829 14656 8893 14660
rect 8909 14716 8973 14720
rect 8909 14660 8913 14716
rect 8913 14660 8969 14716
rect 8969 14660 8973 14716
rect 8909 14656 8973 14660
rect 8989 14716 9053 14720
rect 8989 14660 8993 14716
rect 8993 14660 9049 14716
rect 9049 14660 9053 14716
rect 8989 14656 9053 14660
rect 9069 14716 9133 14720
rect 9069 14660 9073 14716
rect 9073 14660 9129 14716
rect 9129 14660 9133 14716
rect 9069 14656 9133 14660
rect 11980 14716 12044 14720
rect 11980 14660 11984 14716
rect 11984 14660 12040 14716
rect 12040 14660 12044 14716
rect 11980 14656 12044 14660
rect 12060 14716 12124 14720
rect 12060 14660 12064 14716
rect 12064 14660 12120 14716
rect 12120 14660 12124 14716
rect 12060 14656 12124 14660
rect 12140 14716 12204 14720
rect 12140 14660 12144 14716
rect 12144 14660 12200 14716
rect 12200 14660 12204 14716
rect 12140 14656 12204 14660
rect 12220 14716 12284 14720
rect 12220 14660 12224 14716
rect 12224 14660 12280 14716
rect 12280 14660 12284 14716
rect 12220 14656 12284 14660
rect 3187 14172 3251 14176
rect 3187 14116 3191 14172
rect 3191 14116 3247 14172
rect 3247 14116 3251 14172
rect 3187 14112 3251 14116
rect 3267 14172 3331 14176
rect 3267 14116 3271 14172
rect 3271 14116 3327 14172
rect 3327 14116 3331 14172
rect 3267 14112 3331 14116
rect 3347 14172 3411 14176
rect 3347 14116 3351 14172
rect 3351 14116 3407 14172
rect 3407 14116 3411 14172
rect 3347 14112 3411 14116
rect 3427 14172 3491 14176
rect 3427 14116 3431 14172
rect 3431 14116 3487 14172
rect 3487 14116 3491 14172
rect 3427 14112 3491 14116
rect 6338 14172 6402 14176
rect 6338 14116 6342 14172
rect 6342 14116 6398 14172
rect 6398 14116 6402 14172
rect 6338 14112 6402 14116
rect 6418 14172 6482 14176
rect 6418 14116 6422 14172
rect 6422 14116 6478 14172
rect 6478 14116 6482 14172
rect 6418 14112 6482 14116
rect 6498 14172 6562 14176
rect 6498 14116 6502 14172
rect 6502 14116 6558 14172
rect 6558 14116 6562 14172
rect 6498 14112 6562 14116
rect 6578 14172 6642 14176
rect 6578 14116 6582 14172
rect 6582 14116 6638 14172
rect 6638 14116 6642 14172
rect 6578 14112 6642 14116
rect 9489 14172 9553 14176
rect 9489 14116 9493 14172
rect 9493 14116 9549 14172
rect 9549 14116 9553 14172
rect 9489 14112 9553 14116
rect 9569 14172 9633 14176
rect 9569 14116 9573 14172
rect 9573 14116 9629 14172
rect 9629 14116 9633 14172
rect 9569 14112 9633 14116
rect 9649 14172 9713 14176
rect 9649 14116 9653 14172
rect 9653 14116 9709 14172
rect 9709 14116 9713 14172
rect 9649 14112 9713 14116
rect 9729 14172 9793 14176
rect 9729 14116 9733 14172
rect 9733 14116 9789 14172
rect 9789 14116 9793 14172
rect 9729 14112 9793 14116
rect 12640 14172 12704 14176
rect 12640 14116 12644 14172
rect 12644 14116 12700 14172
rect 12700 14116 12704 14172
rect 12640 14112 12704 14116
rect 12720 14172 12784 14176
rect 12720 14116 12724 14172
rect 12724 14116 12780 14172
rect 12780 14116 12784 14172
rect 12720 14112 12784 14116
rect 12800 14172 12864 14176
rect 12800 14116 12804 14172
rect 12804 14116 12860 14172
rect 12860 14116 12864 14172
rect 12800 14112 12864 14116
rect 12880 14172 12944 14176
rect 12880 14116 12884 14172
rect 12884 14116 12940 14172
rect 12940 14116 12944 14172
rect 12880 14112 12944 14116
rect 2527 13628 2591 13632
rect 2527 13572 2531 13628
rect 2531 13572 2587 13628
rect 2587 13572 2591 13628
rect 2527 13568 2591 13572
rect 2607 13628 2671 13632
rect 2607 13572 2611 13628
rect 2611 13572 2667 13628
rect 2667 13572 2671 13628
rect 2607 13568 2671 13572
rect 2687 13628 2751 13632
rect 2687 13572 2691 13628
rect 2691 13572 2747 13628
rect 2747 13572 2751 13628
rect 2687 13568 2751 13572
rect 2767 13628 2831 13632
rect 2767 13572 2771 13628
rect 2771 13572 2827 13628
rect 2827 13572 2831 13628
rect 2767 13568 2831 13572
rect 5678 13628 5742 13632
rect 5678 13572 5682 13628
rect 5682 13572 5738 13628
rect 5738 13572 5742 13628
rect 5678 13568 5742 13572
rect 5758 13628 5822 13632
rect 5758 13572 5762 13628
rect 5762 13572 5818 13628
rect 5818 13572 5822 13628
rect 5758 13568 5822 13572
rect 5838 13628 5902 13632
rect 5838 13572 5842 13628
rect 5842 13572 5898 13628
rect 5898 13572 5902 13628
rect 5838 13568 5902 13572
rect 5918 13628 5982 13632
rect 5918 13572 5922 13628
rect 5922 13572 5978 13628
rect 5978 13572 5982 13628
rect 5918 13568 5982 13572
rect 8829 13628 8893 13632
rect 8829 13572 8833 13628
rect 8833 13572 8889 13628
rect 8889 13572 8893 13628
rect 8829 13568 8893 13572
rect 8909 13628 8973 13632
rect 8909 13572 8913 13628
rect 8913 13572 8969 13628
rect 8969 13572 8973 13628
rect 8909 13568 8973 13572
rect 8989 13628 9053 13632
rect 8989 13572 8993 13628
rect 8993 13572 9049 13628
rect 9049 13572 9053 13628
rect 8989 13568 9053 13572
rect 9069 13628 9133 13632
rect 9069 13572 9073 13628
rect 9073 13572 9129 13628
rect 9129 13572 9133 13628
rect 9069 13568 9133 13572
rect 11980 13628 12044 13632
rect 11980 13572 11984 13628
rect 11984 13572 12040 13628
rect 12040 13572 12044 13628
rect 11980 13568 12044 13572
rect 12060 13628 12124 13632
rect 12060 13572 12064 13628
rect 12064 13572 12120 13628
rect 12120 13572 12124 13628
rect 12060 13568 12124 13572
rect 12140 13628 12204 13632
rect 12140 13572 12144 13628
rect 12144 13572 12200 13628
rect 12200 13572 12204 13628
rect 12140 13568 12204 13572
rect 12220 13628 12284 13632
rect 12220 13572 12224 13628
rect 12224 13572 12280 13628
rect 12280 13572 12284 13628
rect 12220 13568 12284 13572
rect 3187 13084 3251 13088
rect 3187 13028 3191 13084
rect 3191 13028 3247 13084
rect 3247 13028 3251 13084
rect 3187 13024 3251 13028
rect 3267 13084 3331 13088
rect 3267 13028 3271 13084
rect 3271 13028 3327 13084
rect 3327 13028 3331 13084
rect 3267 13024 3331 13028
rect 3347 13084 3411 13088
rect 3347 13028 3351 13084
rect 3351 13028 3407 13084
rect 3407 13028 3411 13084
rect 3347 13024 3411 13028
rect 3427 13084 3491 13088
rect 3427 13028 3431 13084
rect 3431 13028 3487 13084
rect 3487 13028 3491 13084
rect 3427 13024 3491 13028
rect 6338 13084 6402 13088
rect 6338 13028 6342 13084
rect 6342 13028 6398 13084
rect 6398 13028 6402 13084
rect 6338 13024 6402 13028
rect 6418 13084 6482 13088
rect 6418 13028 6422 13084
rect 6422 13028 6478 13084
rect 6478 13028 6482 13084
rect 6418 13024 6482 13028
rect 6498 13084 6562 13088
rect 6498 13028 6502 13084
rect 6502 13028 6558 13084
rect 6558 13028 6562 13084
rect 6498 13024 6562 13028
rect 6578 13084 6642 13088
rect 6578 13028 6582 13084
rect 6582 13028 6638 13084
rect 6638 13028 6642 13084
rect 6578 13024 6642 13028
rect 9489 13084 9553 13088
rect 9489 13028 9493 13084
rect 9493 13028 9549 13084
rect 9549 13028 9553 13084
rect 9489 13024 9553 13028
rect 9569 13084 9633 13088
rect 9569 13028 9573 13084
rect 9573 13028 9629 13084
rect 9629 13028 9633 13084
rect 9569 13024 9633 13028
rect 9649 13084 9713 13088
rect 9649 13028 9653 13084
rect 9653 13028 9709 13084
rect 9709 13028 9713 13084
rect 9649 13024 9713 13028
rect 9729 13084 9793 13088
rect 9729 13028 9733 13084
rect 9733 13028 9789 13084
rect 9789 13028 9793 13084
rect 9729 13024 9793 13028
rect 12640 13084 12704 13088
rect 12640 13028 12644 13084
rect 12644 13028 12700 13084
rect 12700 13028 12704 13084
rect 12640 13024 12704 13028
rect 12720 13084 12784 13088
rect 12720 13028 12724 13084
rect 12724 13028 12780 13084
rect 12780 13028 12784 13084
rect 12720 13024 12784 13028
rect 12800 13084 12864 13088
rect 12800 13028 12804 13084
rect 12804 13028 12860 13084
rect 12860 13028 12864 13084
rect 12800 13024 12864 13028
rect 12880 13084 12944 13088
rect 12880 13028 12884 13084
rect 12884 13028 12940 13084
rect 12940 13028 12944 13084
rect 12880 13024 12944 13028
rect 2527 12540 2591 12544
rect 2527 12484 2531 12540
rect 2531 12484 2587 12540
rect 2587 12484 2591 12540
rect 2527 12480 2591 12484
rect 2607 12540 2671 12544
rect 2607 12484 2611 12540
rect 2611 12484 2667 12540
rect 2667 12484 2671 12540
rect 2607 12480 2671 12484
rect 2687 12540 2751 12544
rect 2687 12484 2691 12540
rect 2691 12484 2747 12540
rect 2747 12484 2751 12540
rect 2687 12480 2751 12484
rect 2767 12540 2831 12544
rect 2767 12484 2771 12540
rect 2771 12484 2827 12540
rect 2827 12484 2831 12540
rect 2767 12480 2831 12484
rect 5678 12540 5742 12544
rect 5678 12484 5682 12540
rect 5682 12484 5738 12540
rect 5738 12484 5742 12540
rect 5678 12480 5742 12484
rect 5758 12540 5822 12544
rect 5758 12484 5762 12540
rect 5762 12484 5818 12540
rect 5818 12484 5822 12540
rect 5758 12480 5822 12484
rect 5838 12540 5902 12544
rect 5838 12484 5842 12540
rect 5842 12484 5898 12540
rect 5898 12484 5902 12540
rect 5838 12480 5902 12484
rect 5918 12540 5982 12544
rect 5918 12484 5922 12540
rect 5922 12484 5978 12540
rect 5978 12484 5982 12540
rect 5918 12480 5982 12484
rect 8829 12540 8893 12544
rect 8829 12484 8833 12540
rect 8833 12484 8889 12540
rect 8889 12484 8893 12540
rect 8829 12480 8893 12484
rect 8909 12540 8973 12544
rect 8909 12484 8913 12540
rect 8913 12484 8969 12540
rect 8969 12484 8973 12540
rect 8909 12480 8973 12484
rect 8989 12540 9053 12544
rect 8989 12484 8993 12540
rect 8993 12484 9049 12540
rect 9049 12484 9053 12540
rect 8989 12480 9053 12484
rect 9069 12540 9133 12544
rect 9069 12484 9073 12540
rect 9073 12484 9129 12540
rect 9129 12484 9133 12540
rect 9069 12480 9133 12484
rect 11980 12540 12044 12544
rect 11980 12484 11984 12540
rect 11984 12484 12040 12540
rect 12040 12484 12044 12540
rect 11980 12480 12044 12484
rect 12060 12540 12124 12544
rect 12060 12484 12064 12540
rect 12064 12484 12120 12540
rect 12120 12484 12124 12540
rect 12060 12480 12124 12484
rect 12140 12540 12204 12544
rect 12140 12484 12144 12540
rect 12144 12484 12200 12540
rect 12200 12484 12204 12540
rect 12140 12480 12204 12484
rect 12220 12540 12284 12544
rect 12220 12484 12224 12540
rect 12224 12484 12280 12540
rect 12280 12484 12284 12540
rect 12220 12480 12284 12484
rect 6132 12276 6196 12340
rect 3187 11996 3251 12000
rect 3187 11940 3191 11996
rect 3191 11940 3247 11996
rect 3247 11940 3251 11996
rect 3187 11936 3251 11940
rect 3267 11996 3331 12000
rect 3267 11940 3271 11996
rect 3271 11940 3327 11996
rect 3327 11940 3331 11996
rect 3267 11936 3331 11940
rect 3347 11996 3411 12000
rect 3347 11940 3351 11996
rect 3351 11940 3407 11996
rect 3407 11940 3411 11996
rect 3347 11936 3411 11940
rect 3427 11996 3491 12000
rect 3427 11940 3431 11996
rect 3431 11940 3487 11996
rect 3487 11940 3491 11996
rect 3427 11936 3491 11940
rect 6338 11996 6402 12000
rect 6338 11940 6342 11996
rect 6342 11940 6398 11996
rect 6398 11940 6402 11996
rect 6338 11936 6402 11940
rect 6418 11996 6482 12000
rect 6418 11940 6422 11996
rect 6422 11940 6478 11996
rect 6478 11940 6482 11996
rect 6418 11936 6482 11940
rect 6498 11996 6562 12000
rect 6498 11940 6502 11996
rect 6502 11940 6558 11996
rect 6558 11940 6562 11996
rect 6498 11936 6562 11940
rect 6578 11996 6642 12000
rect 6578 11940 6582 11996
rect 6582 11940 6638 11996
rect 6638 11940 6642 11996
rect 6578 11936 6642 11940
rect 9489 11996 9553 12000
rect 9489 11940 9493 11996
rect 9493 11940 9549 11996
rect 9549 11940 9553 11996
rect 9489 11936 9553 11940
rect 9569 11996 9633 12000
rect 9569 11940 9573 11996
rect 9573 11940 9629 11996
rect 9629 11940 9633 11996
rect 9569 11936 9633 11940
rect 9649 11996 9713 12000
rect 9649 11940 9653 11996
rect 9653 11940 9709 11996
rect 9709 11940 9713 11996
rect 9649 11936 9713 11940
rect 9729 11996 9793 12000
rect 9729 11940 9733 11996
rect 9733 11940 9789 11996
rect 9789 11940 9793 11996
rect 9729 11936 9793 11940
rect 12640 11996 12704 12000
rect 12640 11940 12644 11996
rect 12644 11940 12700 11996
rect 12700 11940 12704 11996
rect 12640 11936 12704 11940
rect 12720 11996 12784 12000
rect 12720 11940 12724 11996
rect 12724 11940 12780 11996
rect 12780 11940 12784 11996
rect 12720 11936 12784 11940
rect 12800 11996 12864 12000
rect 12800 11940 12804 11996
rect 12804 11940 12860 11996
rect 12860 11940 12864 11996
rect 12800 11936 12864 11940
rect 12880 11996 12944 12000
rect 12880 11940 12884 11996
rect 12884 11940 12940 11996
rect 12940 11940 12944 11996
rect 12880 11936 12944 11940
rect 2527 11452 2591 11456
rect 2527 11396 2531 11452
rect 2531 11396 2587 11452
rect 2587 11396 2591 11452
rect 2527 11392 2591 11396
rect 2607 11452 2671 11456
rect 2607 11396 2611 11452
rect 2611 11396 2667 11452
rect 2667 11396 2671 11452
rect 2607 11392 2671 11396
rect 2687 11452 2751 11456
rect 2687 11396 2691 11452
rect 2691 11396 2747 11452
rect 2747 11396 2751 11452
rect 2687 11392 2751 11396
rect 2767 11452 2831 11456
rect 2767 11396 2771 11452
rect 2771 11396 2827 11452
rect 2827 11396 2831 11452
rect 2767 11392 2831 11396
rect 5678 11452 5742 11456
rect 5678 11396 5682 11452
rect 5682 11396 5738 11452
rect 5738 11396 5742 11452
rect 5678 11392 5742 11396
rect 5758 11452 5822 11456
rect 5758 11396 5762 11452
rect 5762 11396 5818 11452
rect 5818 11396 5822 11452
rect 5758 11392 5822 11396
rect 5838 11452 5902 11456
rect 5838 11396 5842 11452
rect 5842 11396 5898 11452
rect 5898 11396 5902 11452
rect 5838 11392 5902 11396
rect 5918 11452 5982 11456
rect 5918 11396 5922 11452
rect 5922 11396 5978 11452
rect 5978 11396 5982 11452
rect 5918 11392 5982 11396
rect 8829 11452 8893 11456
rect 8829 11396 8833 11452
rect 8833 11396 8889 11452
rect 8889 11396 8893 11452
rect 8829 11392 8893 11396
rect 8909 11452 8973 11456
rect 8909 11396 8913 11452
rect 8913 11396 8969 11452
rect 8969 11396 8973 11452
rect 8909 11392 8973 11396
rect 8989 11452 9053 11456
rect 8989 11396 8993 11452
rect 8993 11396 9049 11452
rect 9049 11396 9053 11452
rect 8989 11392 9053 11396
rect 9069 11452 9133 11456
rect 9069 11396 9073 11452
rect 9073 11396 9129 11452
rect 9129 11396 9133 11452
rect 9069 11392 9133 11396
rect 11980 11452 12044 11456
rect 11980 11396 11984 11452
rect 11984 11396 12040 11452
rect 12040 11396 12044 11452
rect 11980 11392 12044 11396
rect 12060 11452 12124 11456
rect 12060 11396 12064 11452
rect 12064 11396 12120 11452
rect 12120 11396 12124 11452
rect 12060 11392 12124 11396
rect 12140 11452 12204 11456
rect 12140 11396 12144 11452
rect 12144 11396 12200 11452
rect 12200 11396 12204 11452
rect 12140 11392 12204 11396
rect 12220 11452 12284 11456
rect 12220 11396 12224 11452
rect 12224 11396 12280 11452
rect 12280 11396 12284 11452
rect 12220 11392 12284 11396
rect 3187 10908 3251 10912
rect 3187 10852 3191 10908
rect 3191 10852 3247 10908
rect 3247 10852 3251 10908
rect 3187 10848 3251 10852
rect 3267 10908 3331 10912
rect 3267 10852 3271 10908
rect 3271 10852 3327 10908
rect 3327 10852 3331 10908
rect 3267 10848 3331 10852
rect 3347 10908 3411 10912
rect 3347 10852 3351 10908
rect 3351 10852 3407 10908
rect 3407 10852 3411 10908
rect 3347 10848 3411 10852
rect 3427 10908 3491 10912
rect 3427 10852 3431 10908
rect 3431 10852 3487 10908
rect 3487 10852 3491 10908
rect 3427 10848 3491 10852
rect 6338 10908 6402 10912
rect 6338 10852 6342 10908
rect 6342 10852 6398 10908
rect 6398 10852 6402 10908
rect 6338 10848 6402 10852
rect 6418 10908 6482 10912
rect 6418 10852 6422 10908
rect 6422 10852 6478 10908
rect 6478 10852 6482 10908
rect 6418 10848 6482 10852
rect 6498 10908 6562 10912
rect 6498 10852 6502 10908
rect 6502 10852 6558 10908
rect 6558 10852 6562 10908
rect 6498 10848 6562 10852
rect 6578 10908 6642 10912
rect 6578 10852 6582 10908
rect 6582 10852 6638 10908
rect 6638 10852 6642 10908
rect 6578 10848 6642 10852
rect 9489 10908 9553 10912
rect 9489 10852 9493 10908
rect 9493 10852 9549 10908
rect 9549 10852 9553 10908
rect 9489 10848 9553 10852
rect 9569 10908 9633 10912
rect 9569 10852 9573 10908
rect 9573 10852 9629 10908
rect 9629 10852 9633 10908
rect 9569 10848 9633 10852
rect 9649 10908 9713 10912
rect 9649 10852 9653 10908
rect 9653 10852 9709 10908
rect 9709 10852 9713 10908
rect 9649 10848 9713 10852
rect 9729 10908 9793 10912
rect 9729 10852 9733 10908
rect 9733 10852 9789 10908
rect 9789 10852 9793 10908
rect 9729 10848 9793 10852
rect 12640 10908 12704 10912
rect 12640 10852 12644 10908
rect 12644 10852 12700 10908
rect 12700 10852 12704 10908
rect 12640 10848 12704 10852
rect 12720 10908 12784 10912
rect 12720 10852 12724 10908
rect 12724 10852 12780 10908
rect 12780 10852 12784 10908
rect 12720 10848 12784 10852
rect 12800 10908 12864 10912
rect 12800 10852 12804 10908
rect 12804 10852 12860 10908
rect 12860 10852 12864 10908
rect 12800 10848 12864 10852
rect 12880 10908 12944 10912
rect 12880 10852 12884 10908
rect 12884 10852 12940 10908
rect 12940 10852 12944 10908
rect 12880 10848 12944 10852
rect 2527 10364 2591 10368
rect 2527 10308 2531 10364
rect 2531 10308 2587 10364
rect 2587 10308 2591 10364
rect 2527 10304 2591 10308
rect 2607 10364 2671 10368
rect 2607 10308 2611 10364
rect 2611 10308 2667 10364
rect 2667 10308 2671 10364
rect 2607 10304 2671 10308
rect 2687 10364 2751 10368
rect 2687 10308 2691 10364
rect 2691 10308 2747 10364
rect 2747 10308 2751 10364
rect 2687 10304 2751 10308
rect 2767 10364 2831 10368
rect 2767 10308 2771 10364
rect 2771 10308 2827 10364
rect 2827 10308 2831 10364
rect 2767 10304 2831 10308
rect 5678 10364 5742 10368
rect 5678 10308 5682 10364
rect 5682 10308 5738 10364
rect 5738 10308 5742 10364
rect 5678 10304 5742 10308
rect 5758 10364 5822 10368
rect 5758 10308 5762 10364
rect 5762 10308 5818 10364
rect 5818 10308 5822 10364
rect 5758 10304 5822 10308
rect 5838 10364 5902 10368
rect 5838 10308 5842 10364
rect 5842 10308 5898 10364
rect 5898 10308 5902 10364
rect 5838 10304 5902 10308
rect 5918 10364 5982 10368
rect 5918 10308 5922 10364
rect 5922 10308 5978 10364
rect 5978 10308 5982 10364
rect 5918 10304 5982 10308
rect 8829 10364 8893 10368
rect 8829 10308 8833 10364
rect 8833 10308 8889 10364
rect 8889 10308 8893 10364
rect 8829 10304 8893 10308
rect 8909 10364 8973 10368
rect 8909 10308 8913 10364
rect 8913 10308 8969 10364
rect 8969 10308 8973 10364
rect 8909 10304 8973 10308
rect 8989 10364 9053 10368
rect 8989 10308 8993 10364
rect 8993 10308 9049 10364
rect 9049 10308 9053 10364
rect 8989 10304 9053 10308
rect 9069 10364 9133 10368
rect 9069 10308 9073 10364
rect 9073 10308 9129 10364
rect 9129 10308 9133 10364
rect 9069 10304 9133 10308
rect 11980 10364 12044 10368
rect 11980 10308 11984 10364
rect 11984 10308 12040 10364
rect 12040 10308 12044 10364
rect 11980 10304 12044 10308
rect 12060 10364 12124 10368
rect 12060 10308 12064 10364
rect 12064 10308 12120 10364
rect 12120 10308 12124 10364
rect 12060 10304 12124 10308
rect 12140 10364 12204 10368
rect 12140 10308 12144 10364
rect 12144 10308 12200 10364
rect 12200 10308 12204 10364
rect 12140 10304 12204 10308
rect 12220 10364 12284 10368
rect 12220 10308 12224 10364
rect 12224 10308 12280 10364
rect 12280 10308 12284 10364
rect 12220 10304 12284 10308
rect 3187 9820 3251 9824
rect 3187 9764 3191 9820
rect 3191 9764 3247 9820
rect 3247 9764 3251 9820
rect 3187 9760 3251 9764
rect 3267 9820 3331 9824
rect 3267 9764 3271 9820
rect 3271 9764 3327 9820
rect 3327 9764 3331 9820
rect 3267 9760 3331 9764
rect 3347 9820 3411 9824
rect 3347 9764 3351 9820
rect 3351 9764 3407 9820
rect 3407 9764 3411 9820
rect 3347 9760 3411 9764
rect 3427 9820 3491 9824
rect 3427 9764 3431 9820
rect 3431 9764 3487 9820
rect 3487 9764 3491 9820
rect 3427 9760 3491 9764
rect 6338 9820 6402 9824
rect 6338 9764 6342 9820
rect 6342 9764 6398 9820
rect 6398 9764 6402 9820
rect 6338 9760 6402 9764
rect 6418 9820 6482 9824
rect 6418 9764 6422 9820
rect 6422 9764 6478 9820
rect 6478 9764 6482 9820
rect 6418 9760 6482 9764
rect 6498 9820 6562 9824
rect 6498 9764 6502 9820
rect 6502 9764 6558 9820
rect 6558 9764 6562 9820
rect 6498 9760 6562 9764
rect 6578 9820 6642 9824
rect 6578 9764 6582 9820
rect 6582 9764 6638 9820
rect 6638 9764 6642 9820
rect 6578 9760 6642 9764
rect 9489 9820 9553 9824
rect 9489 9764 9493 9820
rect 9493 9764 9549 9820
rect 9549 9764 9553 9820
rect 9489 9760 9553 9764
rect 9569 9820 9633 9824
rect 9569 9764 9573 9820
rect 9573 9764 9629 9820
rect 9629 9764 9633 9820
rect 9569 9760 9633 9764
rect 9649 9820 9713 9824
rect 9649 9764 9653 9820
rect 9653 9764 9709 9820
rect 9709 9764 9713 9820
rect 9649 9760 9713 9764
rect 9729 9820 9793 9824
rect 9729 9764 9733 9820
rect 9733 9764 9789 9820
rect 9789 9764 9793 9820
rect 9729 9760 9793 9764
rect 12640 9820 12704 9824
rect 12640 9764 12644 9820
rect 12644 9764 12700 9820
rect 12700 9764 12704 9820
rect 12640 9760 12704 9764
rect 12720 9820 12784 9824
rect 12720 9764 12724 9820
rect 12724 9764 12780 9820
rect 12780 9764 12784 9820
rect 12720 9760 12784 9764
rect 12800 9820 12864 9824
rect 12800 9764 12804 9820
rect 12804 9764 12860 9820
rect 12860 9764 12864 9820
rect 12800 9760 12864 9764
rect 12880 9820 12944 9824
rect 12880 9764 12884 9820
rect 12884 9764 12940 9820
rect 12940 9764 12944 9820
rect 12880 9760 12944 9764
rect 6132 9556 6196 9620
rect 2527 9276 2591 9280
rect 2527 9220 2531 9276
rect 2531 9220 2587 9276
rect 2587 9220 2591 9276
rect 2527 9216 2591 9220
rect 2607 9276 2671 9280
rect 2607 9220 2611 9276
rect 2611 9220 2667 9276
rect 2667 9220 2671 9276
rect 2607 9216 2671 9220
rect 2687 9276 2751 9280
rect 2687 9220 2691 9276
rect 2691 9220 2747 9276
rect 2747 9220 2751 9276
rect 2687 9216 2751 9220
rect 2767 9276 2831 9280
rect 2767 9220 2771 9276
rect 2771 9220 2827 9276
rect 2827 9220 2831 9276
rect 2767 9216 2831 9220
rect 5678 9276 5742 9280
rect 5678 9220 5682 9276
rect 5682 9220 5738 9276
rect 5738 9220 5742 9276
rect 5678 9216 5742 9220
rect 5758 9276 5822 9280
rect 5758 9220 5762 9276
rect 5762 9220 5818 9276
rect 5818 9220 5822 9276
rect 5758 9216 5822 9220
rect 5838 9276 5902 9280
rect 5838 9220 5842 9276
rect 5842 9220 5898 9276
rect 5898 9220 5902 9276
rect 5838 9216 5902 9220
rect 5918 9276 5982 9280
rect 5918 9220 5922 9276
rect 5922 9220 5978 9276
rect 5978 9220 5982 9276
rect 5918 9216 5982 9220
rect 8829 9276 8893 9280
rect 8829 9220 8833 9276
rect 8833 9220 8889 9276
rect 8889 9220 8893 9276
rect 8829 9216 8893 9220
rect 8909 9276 8973 9280
rect 8909 9220 8913 9276
rect 8913 9220 8969 9276
rect 8969 9220 8973 9276
rect 8909 9216 8973 9220
rect 8989 9276 9053 9280
rect 8989 9220 8993 9276
rect 8993 9220 9049 9276
rect 9049 9220 9053 9276
rect 8989 9216 9053 9220
rect 9069 9276 9133 9280
rect 9069 9220 9073 9276
rect 9073 9220 9129 9276
rect 9129 9220 9133 9276
rect 9069 9216 9133 9220
rect 11980 9276 12044 9280
rect 11980 9220 11984 9276
rect 11984 9220 12040 9276
rect 12040 9220 12044 9276
rect 11980 9216 12044 9220
rect 12060 9276 12124 9280
rect 12060 9220 12064 9276
rect 12064 9220 12120 9276
rect 12120 9220 12124 9276
rect 12060 9216 12124 9220
rect 12140 9276 12204 9280
rect 12140 9220 12144 9276
rect 12144 9220 12200 9276
rect 12200 9220 12204 9276
rect 12140 9216 12204 9220
rect 12220 9276 12284 9280
rect 12220 9220 12224 9276
rect 12224 9220 12280 9276
rect 12280 9220 12284 9276
rect 12220 9216 12284 9220
rect 3187 8732 3251 8736
rect 3187 8676 3191 8732
rect 3191 8676 3247 8732
rect 3247 8676 3251 8732
rect 3187 8672 3251 8676
rect 3267 8732 3331 8736
rect 3267 8676 3271 8732
rect 3271 8676 3327 8732
rect 3327 8676 3331 8732
rect 3267 8672 3331 8676
rect 3347 8732 3411 8736
rect 3347 8676 3351 8732
rect 3351 8676 3407 8732
rect 3407 8676 3411 8732
rect 3347 8672 3411 8676
rect 3427 8732 3491 8736
rect 3427 8676 3431 8732
rect 3431 8676 3487 8732
rect 3487 8676 3491 8732
rect 3427 8672 3491 8676
rect 6338 8732 6402 8736
rect 6338 8676 6342 8732
rect 6342 8676 6398 8732
rect 6398 8676 6402 8732
rect 6338 8672 6402 8676
rect 6418 8732 6482 8736
rect 6418 8676 6422 8732
rect 6422 8676 6478 8732
rect 6478 8676 6482 8732
rect 6418 8672 6482 8676
rect 6498 8732 6562 8736
rect 6498 8676 6502 8732
rect 6502 8676 6558 8732
rect 6558 8676 6562 8732
rect 6498 8672 6562 8676
rect 6578 8732 6642 8736
rect 6578 8676 6582 8732
rect 6582 8676 6638 8732
rect 6638 8676 6642 8732
rect 6578 8672 6642 8676
rect 9489 8732 9553 8736
rect 9489 8676 9493 8732
rect 9493 8676 9549 8732
rect 9549 8676 9553 8732
rect 9489 8672 9553 8676
rect 9569 8732 9633 8736
rect 9569 8676 9573 8732
rect 9573 8676 9629 8732
rect 9629 8676 9633 8732
rect 9569 8672 9633 8676
rect 9649 8732 9713 8736
rect 9649 8676 9653 8732
rect 9653 8676 9709 8732
rect 9709 8676 9713 8732
rect 9649 8672 9713 8676
rect 9729 8732 9793 8736
rect 9729 8676 9733 8732
rect 9733 8676 9789 8732
rect 9789 8676 9793 8732
rect 9729 8672 9793 8676
rect 12640 8732 12704 8736
rect 12640 8676 12644 8732
rect 12644 8676 12700 8732
rect 12700 8676 12704 8732
rect 12640 8672 12704 8676
rect 12720 8732 12784 8736
rect 12720 8676 12724 8732
rect 12724 8676 12780 8732
rect 12780 8676 12784 8732
rect 12720 8672 12784 8676
rect 12800 8732 12864 8736
rect 12800 8676 12804 8732
rect 12804 8676 12860 8732
rect 12860 8676 12864 8732
rect 12800 8672 12864 8676
rect 12880 8732 12944 8736
rect 12880 8676 12884 8732
rect 12884 8676 12940 8732
rect 12940 8676 12944 8732
rect 12880 8672 12944 8676
rect 2527 8188 2591 8192
rect 2527 8132 2531 8188
rect 2531 8132 2587 8188
rect 2587 8132 2591 8188
rect 2527 8128 2591 8132
rect 2607 8188 2671 8192
rect 2607 8132 2611 8188
rect 2611 8132 2667 8188
rect 2667 8132 2671 8188
rect 2607 8128 2671 8132
rect 2687 8188 2751 8192
rect 2687 8132 2691 8188
rect 2691 8132 2747 8188
rect 2747 8132 2751 8188
rect 2687 8128 2751 8132
rect 2767 8188 2831 8192
rect 2767 8132 2771 8188
rect 2771 8132 2827 8188
rect 2827 8132 2831 8188
rect 2767 8128 2831 8132
rect 5678 8188 5742 8192
rect 5678 8132 5682 8188
rect 5682 8132 5738 8188
rect 5738 8132 5742 8188
rect 5678 8128 5742 8132
rect 5758 8188 5822 8192
rect 5758 8132 5762 8188
rect 5762 8132 5818 8188
rect 5818 8132 5822 8188
rect 5758 8128 5822 8132
rect 5838 8188 5902 8192
rect 5838 8132 5842 8188
rect 5842 8132 5898 8188
rect 5898 8132 5902 8188
rect 5838 8128 5902 8132
rect 5918 8188 5982 8192
rect 5918 8132 5922 8188
rect 5922 8132 5978 8188
rect 5978 8132 5982 8188
rect 5918 8128 5982 8132
rect 8829 8188 8893 8192
rect 8829 8132 8833 8188
rect 8833 8132 8889 8188
rect 8889 8132 8893 8188
rect 8829 8128 8893 8132
rect 8909 8188 8973 8192
rect 8909 8132 8913 8188
rect 8913 8132 8969 8188
rect 8969 8132 8973 8188
rect 8909 8128 8973 8132
rect 8989 8188 9053 8192
rect 8989 8132 8993 8188
rect 8993 8132 9049 8188
rect 9049 8132 9053 8188
rect 8989 8128 9053 8132
rect 9069 8188 9133 8192
rect 9069 8132 9073 8188
rect 9073 8132 9129 8188
rect 9129 8132 9133 8188
rect 9069 8128 9133 8132
rect 11980 8188 12044 8192
rect 11980 8132 11984 8188
rect 11984 8132 12040 8188
rect 12040 8132 12044 8188
rect 11980 8128 12044 8132
rect 12060 8188 12124 8192
rect 12060 8132 12064 8188
rect 12064 8132 12120 8188
rect 12120 8132 12124 8188
rect 12060 8128 12124 8132
rect 12140 8188 12204 8192
rect 12140 8132 12144 8188
rect 12144 8132 12200 8188
rect 12200 8132 12204 8188
rect 12140 8128 12204 8132
rect 12220 8188 12284 8192
rect 12220 8132 12224 8188
rect 12224 8132 12280 8188
rect 12280 8132 12284 8188
rect 12220 8128 12284 8132
rect 3187 7644 3251 7648
rect 3187 7588 3191 7644
rect 3191 7588 3247 7644
rect 3247 7588 3251 7644
rect 3187 7584 3251 7588
rect 3267 7644 3331 7648
rect 3267 7588 3271 7644
rect 3271 7588 3327 7644
rect 3327 7588 3331 7644
rect 3267 7584 3331 7588
rect 3347 7644 3411 7648
rect 3347 7588 3351 7644
rect 3351 7588 3407 7644
rect 3407 7588 3411 7644
rect 3347 7584 3411 7588
rect 3427 7644 3491 7648
rect 3427 7588 3431 7644
rect 3431 7588 3487 7644
rect 3487 7588 3491 7644
rect 3427 7584 3491 7588
rect 6338 7644 6402 7648
rect 6338 7588 6342 7644
rect 6342 7588 6398 7644
rect 6398 7588 6402 7644
rect 6338 7584 6402 7588
rect 6418 7644 6482 7648
rect 6418 7588 6422 7644
rect 6422 7588 6478 7644
rect 6478 7588 6482 7644
rect 6418 7584 6482 7588
rect 6498 7644 6562 7648
rect 6498 7588 6502 7644
rect 6502 7588 6558 7644
rect 6558 7588 6562 7644
rect 6498 7584 6562 7588
rect 6578 7644 6642 7648
rect 6578 7588 6582 7644
rect 6582 7588 6638 7644
rect 6638 7588 6642 7644
rect 6578 7584 6642 7588
rect 9489 7644 9553 7648
rect 9489 7588 9493 7644
rect 9493 7588 9549 7644
rect 9549 7588 9553 7644
rect 9489 7584 9553 7588
rect 9569 7644 9633 7648
rect 9569 7588 9573 7644
rect 9573 7588 9629 7644
rect 9629 7588 9633 7644
rect 9569 7584 9633 7588
rect 9649 7644 9713 7648
rect 9649 7588 9653 7644
rect 9653 7588 9709 7644
rect 9709 7588 9713 7644
rect 9649 7584 9713 7588
rect 9729 7644 9793 7648
rect 9729 7588 9733 7644
rect 9733 7588 9789 7644
rect 9789 7588 9793 7644
rect 9729 7584 9793 7588
rect 12640 7644 12704 7648
rect 12640 7588 12644 7644
rect 12644 7588 12700 7644
rect 12700 7588 12704 7644
rect 12640 7584 12704 7588
rect 12720 7644 12784 7648
rect 12720 7588 12724 7644
rect 12724 7588 12780 7644
rect 12780 7588 12784 7644
rect 12720 7584 12784 7588
rect 12800 7644 12864 7648
rect 12800 7588 12804 7644
rect 12804 7588 12860 7644
rect 12860 7588 12864 7644
rect 12800 7584 12864 7588
rect 12880 7644 12944 7648
rect 12880 7588 12884 7644
rect 12884 7588 12940 7644
rect 12940 7588 12944 7644
rect 12880 7584 12944 7588
rect 2527 7100 2591 7104
rect 2527 7044 2531 7100
rect 2531 7044 2587 7100
rect 2587 7044 2591 7100
rect 2527 7040 2591 7044
rect 2607 7100 2671 7104
rect 2607 7044 2611 7100
rect 2611 7044 2667 7100
rect 2667 7044 2671 7100
rect 2607 7040 2671 7044
rect 2687 7100 2751 7104
rect 2687 7044 2691 7100
rect 2691 7044 2747 7100
rect 2747 7044 2751 7100
rect 2687 7040 2751 7044
rect 2767 7100 2831 7104
rect 2767 7044 2771 7100
rect 2771 7044 2827 7100
rect 2827 7044 2831 7100
rect 2767 7040 2831 7044
rect 5678 7100 5742 7104
rect 5678 7044 5682 7100
rect 5682 7044 5738 7100
rect 5738 7044 5742 7100
rect 5678 7040 5742 7044
rect 5758 7100 5822 7104
rect 5758 7044 5762 7100
rect 5762 7044 5818 7100
rect 5818 7044 5822 7100
rect 5758 7040 5822 7044
rect 5838 7100 5902 7104
rect 5838 7044 5842 7100
rect 5842 7044 5898 7100
rect 5898 7044 5902 7100
rect 5838 7040 5902 7044
rect 5918 7100 5982 7104
rect 5918 7044 5922 7100
rect 5922 7044 5978 7100
rect 5978 7044 5982 7100
rect 5918 7040 5982 7044
rect 8829 7100 8893 7104
rect 8829 7044 8833 7100
rect 8833 7044 8889 7100
rect 8889 7044 8893 7100
rect 8829 7040 8893 7044
rect 8909 7100 8973 7104
rect 8909 7044 8913 7100
rect 8913 7044 8969 7100
rect 8969 7044 8973 7100
rect 8909 7040 8973 7044
rect 8989 7100 9053 7104
rect 8989 7044 8993 7100
rect 8993 7044 9049 7100
rect 9049 7044 9053 7100
rect 8989 7040 9053 7044
rect 9069 7100 9133 7104
rect 9069 7044 9073 7100
rect 9073 7044 9129 7100
rect 9129 7044 9133 7100
rect 9069 7040 9133 7044
rect 11980 7100 12044 7104
rect 11980 7044 11984 7100
rect 11984 7044 12040 7100
rect 12040 7044 12044 7100
rect 11980 7040 12044 7044
rect 12060 7100 12124 7104
rect 12060 7044 12064 7100
rect 12064 7044 12120 7100
rect 12120 7044 12124 7100
rect 12060 7040 12124 7044
rect 12140 7100 12204 7104
rect 12140 7044 12144 7100
rect 12144 7044 12200 7100
rect 12200 7044 12204 7100
rect 12140 7040 12204 7044
rect 12220 7100 12284 7104
rect 12220 7044 12224 7100
rect 12224 7044 12280 7100
rect 12280 7044 12284 7100
rect 12220 7040 12284 7044
rect 3187 6556 3251 6560
rect 3187 6500 3191 6556
rect 3191 6500 3247 6556
rect 3247 6500 3251 6556
rect 3187 6496 3251 6500
rect 3267 6556 3331 6560
rect 3267 6500 3271 6556
rect 3271 6500 3327 6556
rect 3327 6500 3331 6556
rect 3267 6496 3331 6500
rect 3347 6556 3411 6560
rect 3347 6500 3351 6556
rect 3351 6500 3407 6556
rect 3407 6500 3411 6556
rect 3347 6496 3411 6500
rect 3427 6556 3491 6560
rect 3427 6500 3431 6556
rect 3431 6500 3487 6556
rect 3487 6500 3491 6556
rect 3427 6496 3491 6500
rect 6338 6556 6402 6560
rect 6338 6500 6342 6556
rect 6342 6500 6398 6556
rect 6398 6500 6402 6556
rect 6338 6496 6402 6500
rect 6418 6556 6482 6560
rect 6418 6500 6422 6556
rect 6422 6500 6478 6556
rect 6478 6500 6482 6556
rect 6418 6496 6482 6500
rect 6498 6556 6562 6560
rect 6498 6500 6502 6556
rect 6502 6500 6558 6556
rect 6558 6500 6562 6556
rect 6498 6496 6562 6500
rect 6578 6556 6642 6560
rect 6578 6500 6582 6556
rect 6582 6500 6638 6556
rect 6638 6500 6642 6556
rect 6578 6496 6642 6500
rect 9489 6556 9553 6560
rect 9489 6500 9493 6556
rect 9493 6500 9549 6556
rect 9549 6500 9553 6556
rect 9489 6496 9553 6500
rect 9569 6556 9633 6560
rect 9569 6500 9573 6556
rect 9573 6500 9629 6556
rect 9629 6500 9633 6556
rect 9569 6496 9633 6500
rect 9649 6556 9713 6560
rect 9649 6500 9653 6556
rect 9653 6500 9709 6556
rect 9709 6500 9713 6556
rect 9649 6496 9713 6500
rect 9729 6556 9793 6560
rect 9729 6500 9733 6556
rect 9733 6500 9789 6556
rect 9789 6500 9793 6556
rect 9729 6496 9793 6500
rect 12640 6556 12704 6560
rect 12640 6500 12644 6556
rect 12644 6500 12700 6556
rect 12700 6500 12704 6556
rect 12640 6496 12704 6500
rect 12720 6556 12784 6560
rect 12720 6500 12724 6556
rect 12724 6500 12780 6556
rect 12780 6500 12784 6556
rect 12720 6496 12784 6500
rect 12800 6556 12864 6560
rect 12800 6500 12804 6556
rect 12804 6500 12860 6556
rect 12860 6500 12864 6556
rect 12800 6496 12864 6500
rect 12880 6556 12944 6560
rect 12880 6500 12884 6556
rect 12884 6500 12940 6556
rect 12940 6500 12944 6556
rect 12880 6496 12944 6500
rect 2527 6012 2591 6016
rect 2527 5956 2531 6012
rect 2531 5956 2587 6012
rect 2587 5956 2591 6012
rect 2527 5952 2591 5956
rect 2607 6012 2671 6016
rect 2607 5956 2611 6012
rect 2611 5956 2667 6012
rect 2667 5956 2671 6012
rect 2607 5952 2671 5956
rect 2687 6012 2751 6016
rect 2687 5956 2691 6012
rect 2691 5956 2747 6012
rect 2747 5956 2751 6012
rect 2687 5952 2751 5956
rect 2767 6012 2831 6016
rect 2767 5956 2771 6012
rect 2771 5956 2827 6012
rect 2827 5956 2831 6012
rect 2767 5952 2831 5956
rect 5678 6012 5742 6016
rect 5678 5956 5682 6012
rect 5682 5956 5738 6012
rect 5738 5956 5742 6012
rect 5678 5952 5742 5956
rect 5758 6012 5822 6016
rect 5758 5956 5762 6012
rect 5762 5956 5818 6012
rect 5818 5956 5822 6012
rect 5758 5952 5822 5956
rect 5838 6012 5902 6016
rect 5838 5956 5842 6012
rect 5842 5956 5898 6012
rect 5898 5956 5902 6012
rect 5838 5952 5902 5956
rect 5918 6012 5982 6016
rect 5918 5956 5922 6012
rect 5922 5956 5978 6012
rect 5978 5956 5982 6012
rect 5918 5952 5982 5956
rect 8829 6012 8893 6016
rect 8829 5956 8833 6012
rect 8833 5956 8889 6012
rect 8889 5956 8893 6012
rect 8829 5952 8893 5956
rect 8909 6012 8973 6016
rect 8909 5956 8913 6012
rect 8913 5956 8969 6012
rect 8969 5956 8973 6012
rect 8909 5952 8973 5956
rect 8989 6012 9053 6016
rect 8989 5956 8993 6012
rect 8993 5956 9049 6012
rect 9049 5956 9053 6012
rect 8989 5952 9053 5956
rect 9069 6012 9133 6016
rect 9069 5956 9073 6012
rect 9073 5956 9129 6012
rect 9129 5956 9133 6012
rect 9069 5952 9133 5956
rect 11980 6012 12044 6016
rect 11980 5956 11984 6012
rect 11984 5956 12040 6012
rect 12040 5956 12044 6012
rect 11980 5952 12044 5956
rect 12060 6012 12124 6016
rect 12060 5956 12064 6012
rect 12064 5956 12120 6012
rect 12120 5956 12124 6012
rect 12060 5952 12124 5956
rect 12140 6012 12204 6016
rect 12140 5956 12144 6012
rect 12144 5956 12200 6012
rect 12200 5956 12204 6012
rect 12140 5952 12204 5956
rect 12220 6012 12284 6016
rect 12220 5956 12224 6012
rect 12224 5956 12280 6012
rect 12280 5956 12284 6012
rect 12220 5952 12284 5956
rect 3187 5468 3251 5472
rect 3187 5412 3191 5468
rect 3191 5412 3247 5468
rect 3247 5412 3251 5468
rect 3187 5408 3251 5412
rect 3267 5468 3331 5472
rect 3267 5412 3271 5468
rect 3271 5412 3327 5468
rect 3327 5412 3331 5468
rect 3267 5408 3331 5412
rect 3347 5468 3411 5472
rect 3347 5412 3351 5468
rect 3351 5412 3407 5468
rect 3407 5412 3411 5468
rect 3347 5408 3411 5412
rect 3427 5468 3491 5472
rect 3427 5412 3431 5468
rect 3431 5412 3487 5468
rect 3487 5412 3491 5468
rect 3427 5408 3491 5412
rect 6338 5468 6402 5472
rect 6338 5412 6342 5468
rect 6342 5412 6398 5468
rect 6398 5412 6402 5468
rect 6338 5408 6402 5412
rect 6418 5468 6482 5472
rect 6418 5412 6422 5468
rect 6422 5412 6478 5468
rect 6478 5412 6482 5468
rect 6418 5408 6482 5412
rect 6498 5468 6562 5472
rect 6498 5412 6502 5468
rect 6502 5412 6558 5468
rect 6558 5412 6562 5468
rect 6498 5408 6562 5412
rect 6578 5468 6642 5472
rect 6578 5412 6582 5468
rect 6582 5412 6638 5468
rect 6638 5412 6642 5468
rect 6578 5408 6642 5412
rect 9489 5468 9553 5472
rect 9489 5412 9493 5468
rect 9493 5412 9549 5468
rect 9549 5412 9553 5468
rect 9489 5408 9553 5412
rect 9569 5468 9633 5472
rect 9569 5412 9573 5468
rect 9573 5412 9629 5468
rect 9629 5412 9633 5468
rect 9569 5408 9633 5412
rect 9649 5468 9713 5472
rect 9649 5412 9653 5468
rect 9653 5412 9709 5468
rect 9709 5412 9713 5468
rect 9649 5408 9713 5412
rect 9729 5468 9793 5472
rect 9729 5412 9733 5468
rect 9733 5412 9789 5468
rect 9789 5412 9793 5468
rect 9729 5408 9793 5412
rect 12640 5468 12704 5472
rect 12640 5412 12644 5468
rect 12644 5412 12700 5468
rect 12700 5412 12704 5468
rect 12640 5408 12704 5412
rect 12720 5468 12784 5472
rect 12720 5412 12724 5468
rect 12724 5412 12780 5468
rect 12780 5412 12784 5468
rect 12720 5408 12784 5412
rect 12800 5468 12864 5472
rect 12800 5412 12804 5468
rect 12804 5412 12860 5468
rect 12860 5412 12864 5468
rect 12800 5408 12864 5412
rect 12880 5468 12944 5472
rect 12880 5412 12884 5468
rect 12884 5412 12940 5468
rect 12940 5412 12944 5468
rect 12880 5408 12944 5412
rect 2527 4924 2591 4928
rect 2527 4868 2531 4924
rect 2531 4868 2587 4924
rect 2587 4868 2591 4924
rect 2527 4864 2591 4868
rect 2607 4924 2671 4928
rect 2607 4868 2611 4924
rect 2611 4868 2667 4924
rect 2667 4868 2671 4924
rect 2607 4864 2671 4868
rect 2687 4924 2751 4928
rect 2687 4868 2691 4924
rect 2691 4868 2747 4924
rect 2747 4868 2751 4924
rect 2687 4864 2751 4868
rect 2767 4924 2831 4928
rect 2767 4868 2771 4924
rect 2771 4868 2827 4924
rect 2827 4868 2831 4924
rect 2767 4864 2831 4868
rect 5678 4924 5742 4928
rect 5678 4868 5682 4924
rect 5682 4868 5738 4924
rect 5738 4868 5742 4924
rect 5678 4864 5742 4868
rect 5758 4924 5822 4928
rect 5758 4868 5762 4924
rect 5762 4868 5818 4924
rect 5818 4868 5822 4924
rect 5758 4864 5822 4868
rect 5838 4924 5902 4928
rect 5838 4868 5842 4924
rect 5842 4868 5898 4924
rect 5898 4868 5902 4924
rect 5838 4864 5902 4868
rect 5918 4924 5982 4928
rect 5918 4868 5922 4924
rect 5922 4868 5978 4924
rect 5978 4868 5982 4924
rect 5918 4864 5982 4868
rect 8829 4924 8893 4928
rect 8829 4868 8833 4924
rect 8833 4868 8889 4924
rect 8889 4868 8893 4924
rect 8829 4864 8893 4868
rect 8909 4924 8973 4928
rect 8909 4868 8913 4924
rect 8913 4868 8969 4924
rect 8969 4868 8973 4924
rect 8909 4864 8973 4868
rect 8989 4924 9053 4928
rect 8989 4868 8993 4924
rect 8993 4868 9049 4924
rect 9049 4868 9053 4924
rect 8989 4864 9053 4868
rect 9069 4924 9133 4928
rect 9069 4868 9073 4924
rect 9073 4868 9129 4924
rect 9129 4868 9133 4924
rect 9069 4864 9133 4868
rect 11980 4924 12044 4928
rect 11980 4868 11984 4924
rect 11984 4868 12040 4924
rect 12040 4868 12044 4924
rect 11980 4864 12044 4868
rect 12060 4924 12124 4928
rect 12060 4868 12064 4924
rect 12064 4868 12120 4924
rect 12120 4868 12124 4924
rect 12060 4864 12124 4868
rect 12140 4924 12204 4928
rect 12140 4868 12144 4924
rect 12144 4868 12200 4924
rect 12200 4868 12204 4924
rect 12140 4864 12204 4868
rect 12220 4924 12284 4928
rect 12220 4868 12224 4924
rect 12224 4868 12280 4924
rect 12280 4868 12284 4924
rect 12220 4864 12284 4868
rect 3187 4380 3251 4384
rect 3187 4324 3191 4380
rect 3191 4324 3247 4380
rect 3247 4324 3251 4380
rect 3187 4320 3251 4324
rect 3267 4380 3331 4384
rect 3267 4324 3271 4380
rect 3271 4324 3327 4380
rect 3327 4324 3331 4380
rect 3267 4320 3331 4324
rect 3347 4380 3411 4384
rect 3347 4324 3351 4380
rect 3351 4324 3407 4380
rect 3407 4324 3411 4380
rect 3347 4320 3411 4324
rect 3427 4380 3491 4384
rect 3427 4324 3431 4380
rect 3431 4324 3487 4380
rect 3487 4324 3491 4380
rect 3427 4320 3491 4324
rect 6338 4380 6402 4384
rect 6338 4324 6342 4380
rect 6342 4324 6398 4380
rect 6398 4324 6402 4380
rect 6338 4320 6402 4324
rect 6418 4380 6482 4384
rect 6418 4324 6422 4380
rect 6422 4324 6478 4380
rect 6478 4324 6482 4380
rect 6418 4320 6482 4324
rect 6498 4380 6562 4384
rect 6498 4324 6502 4380
rect 6502 4324 6558 4380
rect 6558 4324 6562 4380
rect 6498 4320 6562 4324
rect 6578 4380 6642 4384
rect 6578 4324 6582 4380
rect 6582 4324 6638 4380
rect 6638 4324 6642 4380
rect 6578 4320 6642 4324
rect 9489 4380 9553 4384
rect 9489 4324 9493 4380
rect 9493 4324 9549 4380
rect 9549 4324 9553 4380
rect 9489 4320 9553 4324
rect 9569 4380 9633 4384
rect 9569 4324 9573 4380
rect 9573 4324 9629 4380
rect 9629 4324 9633 4380
rect 9569 4320 9633 4324
rect 9649 4380 9713 4384
rect 9649 4324 9653 4380
rect 9653 4324 9709 4380
rect 9709 4324 9713 4380
rect 9649 4320 9713 4324
rect 9729 4380 9793 4384
rect 9729 4324 9733 4380
rect 9733 4324 9789 4380
rect 9789 4324 9793 4380
rect 9729 4320 9793 4324
rect 12640 4380 12704 4384
rect 12640 4324 12644 4380
rect 12644 4324 12700 4380
rect 12700 4324 12704 4380
rect 12640 4320 12704 4324
rect 12720 4380 12784 4384
rect 12720 4324 12724 4380
rect 12724 4324 12780 4380
rect 12780 4324 12784 4380
rect 12720 4320 12784 4324
rect 12800 4380 12864 4384
rect 12800 4324 12804 4380
rect 12804 4324 12860 4380
rect 12860 4324 12864 4380
rect 12800 4320 12864 4324
rect 12880 4380 12944 4384
rect 12880 4324 12884 4380
rect 12884 4324 12940 4380
rect 12940 4324 12944 4380
rect 12880 4320 12944 4324
rect 2527 3836 2591 3840
rect 2527 3780 2531 3836
rect 2531 3780 2587 3836
rect 2587 3780 2591 3836
rect 2527 3776 2591 3780
rect 2607 3836 2671 3840
rect 2607 3780 2611 3836
rect 2611 3780 2667 3836
rect 2667 3780 2671 3836
rect 2607 3776 2671 3780
rect 2687 3836 2751 3840
rect 2687 3780 2691 3836
rect 2691 3780 2747 3836
rect 2747 3780 2751 3836
rect 2687 3776 2751 3780
rect 2767 3836 2831 3840
rect 2767 3780 2771 3836
rect 2771 3780 2827 3836
rect 2827 3780 2831 3836
rect 2767 3776 2831 3780
rect 5678 3836 5742 3840
rect 5678 3780 5682 3836
rect 5682 3780 5738 3836
rect 5738 3780 5742 3836
rect 5678 3776 5742 3780
rect 5758 3836 5822 3840
rect 5758 3780 5762 3836
rect 5762 3780 5818 3836
rect 5818 3780 5822 3836
rect 5758 3776 5822 3780
rect 5838 3836 5902 3840
rect 5838 3780 5842 3836
rect 5842 3780 5898 3836
rect 5898 3780 5902 3836
rect 5838 3776 5902 3780
rect 5918 3836 5982 3840
rect 5918 3780 5922 3836
rect 5922 3780 5978 3836
rect 5978 3780 5982 3836
rect 5918 3776 5982 3780
rect 8829 3836 8893 3840
rect 8829 3780 8833 3836
rect 8833 3780 8889 3836
rect 8889 3780 8893 3836
rect 8829 3776 8893 3780
rect 8909 3836 8973 3840
rect 8909 3780 8913 3836
rect 8913 3780 8969 3836
rect 8969 3780 8973 3836
rect 8909 3776 8973 3780
rect 8989 3836 9053 3840
rect 8989 3780 8993 3836
rect 8993 3780 9049 3836
rect 9049 3780 9053 3836
rect 8989 3776 9053 3780
rect 9069 3836 9133 3840
rect 9069 3780 9073 3836
rect 9073 3780 9129 3836
rect 9129 3780 9133 3836
rect 9069 3776 9133 3780
rect 11980 3836 12044 3840
rect 11980 3780 11984 3836
rect 11984 3780 12040 3836
rect 12040 3780 12044 3836
rect 11980 3776 12044 3780
rect 12060 3836 12124 3840
rect 12060 3780 12064 3836
rect 12064 3780 12120 3836
rect 12120 3780 12124 3836
rect 12060 3776 12124 3780
rect 12140 3836 12204 3840
rect 12140 3780 12144 3836
rect 12144 3780 12200 3836
rect 12200 3780 12204 3836
rect 12140 3776 12204 3780
rect 12220 3836 12284 3840
rect 12220 3780 12224 3836
rect 12224 3780 12280 3836
rect 12280 3780 12284 3836
rect 12220 3776 12284 3780
rect 3187 3292 3251 3296
rect 3187 3236 3191 3292
rect 3191 3236 3247 3292
rect 3247 3236 3251 3292
rect 3187 3232 3251 3236
rect 3267 3292 3331 3296
rect 3267 3236 3271 3292
rect 3271 3236 3327 3292
rect 3327 3236 3331 3292
rect 3267 3232 3331 3236
rect 3347 3292 3411 3296
rect 3347 3236 3351 3292
rect 3351 3236 3407 3292
rect 3407 3236 3411 3292
rect 3347 3232 3411 3236
rect 3427 3292 3491 3296
rect 3427 3236 3431 3292
rect 3431 3236 3487 3292
rect 3487 3236 3491 3292
rect 3427 3232 3491 3236
rect 6338 3292 6402 3296
rect 6338 3236 6342 3292
rect 6342 3236 6398 3292
rect 6398 3236 6402 3292
rect 6338 3232 6402 3236
rect 6418 3292 6482 3296
rect 6418 3236 6422 3292
rect 6422 3236 6478 3292
rect 6478 3236 6482 3292
rect 6418 3232 6482 3236
rect 6498 3292 6562 3296
rect 6498 3236 6502 3292
rect 6502 3236 6558 3292
rect 6558 3236 6562 3292
rect 6498 3232 6562 3236
rect 6578 3292 6642 3296
rect 6578 3236 6582 3292
rect 6582 3236 6638 3292
rect 6638 3236 6642 3292
rect 6578 3232 6642 3236
rect 9489 3292 9553 3296
rect 9489 3236 9493 3292
rect 9493 3236 9549 3292
rect 9549 3236 9553 3292
rect 9489 3232 9553 3236
rect 9569 3292 9633 3296
rect 9569 3236 9573 3292
rect 9573 3236 9629 3292
rect 9629 3236 9633 3292
rect 9569 3232 9633 3236
rect 9649 3292 9713 3296
rect 9649 3236 9653 3292
rect 9653 3236 9709 3292
rect 9709 3236 9713 3292
rect 9649 3232 9713 3236
rect 9729 3292 9793 3296
rect 9729 3236 9733 3292
rect 9733 3236 9789 3292
rect 9789 3236 9793 3292
rect 9729 3232 9793 3236
rect 12640 3292 12704 3296
rect 12640 3236 12644 3292
rect 12644 3236 12700 3292
rect 12700 3236 12704 3292
rect 12640 3232 12704 3236
rect 12720 3292 12784 3296
rect 12720 3236 12724 3292
rect 12724 3236 12780 3292
rect 12780 3236 12784 3292
rect 12720 3232 12784 3236
rect 12800 3292 12864 3296
rect 12800 3236 12804 3292
rect 12804 3236 12860 3292
rect 12860 3236 12864 3292
rect 12800 3232 12864 3236
rect 12880 3292 12944 3296
rect 12880 3236 12884 3292
rect 12884 3236 12940 3292
rect 12940 3236 12944 3292
rect 12880 3232 12944 3236
rect 2527 2748 2591 2752
rect 2527 2692 2531 2748
rect 2531 2692 2587 2748
rect 2587 2692 2591 2748
rect 2527 2688 2591 2692
rect 2607 2748 2671 2752
rect 2607 2692 2611 2748
rect 2611 2692 2667 2748
rect 2667 2692 2671 2748
rect 2607 2688 2671 2692
rect 2687 2748 2751 2752
rect 2687 2692 2691 2748
rect 2691 2692 2747 2748
rect 2747 2692 2751 2748
rect 2687 2688 2751 2692
rect 2767 2748 2831 2752
rect 2767 2692 2771 2748
rect 2771 2692 2827 2748
rect 2827 2692 2831 2748
rect 2767 2688 2831 2692
rect 5678 2748 5742 2752
rect 5678 2692 5682 2748
rect 5682 2692 5738 2748
rect 5738 2692 5742 2748
rect 5678 2688 5742 2692
rect 5758 2748 5822 2752
rect 5758 2692 5762 2748
rect 5762 2692 5818 2748
rect 5818 2692 5822 2748
rect 5758 2688 5822 2692
rect 5838 2748 5902 2752
rect 5838 2692 5842 2748
rect 5842 2692 5898 2748
rect 5898 2692 5902 2748
rect 5838 2688 5902 2692
rect 5918 2748 5982 2752
rect 5918 2692 5922 2748
rect 5922 2692 5978 2748
rect 5978 2692 5982 2748
rect 5918 2688 5982 2692
rect 8829 2748 8893 2752
rect 8829 2692 8833 2748
rect 8833 2692 8889 2748
rect 8889 2692 8893 2748
rect 8829 2688 8893 2692
rect 8909 2748 8973 2752
rect 8909 2692 8913 2748
rect 8913 2692 8969 2748
rect 8969 2692 8973 2748
rect 8909 2688 8973 2692
rect 8989 2748 9053 2752
rect 8989 2692 8993 2748
rect 8993 2692 9049 2748
rect 9049 2692 9053 2748
rect 8989 2688 9053 2692
rect 9069 2748 9133 2752
rect 9069 2692 9073 2748
rect 9073 2692 9129 2748
rect 9129 2692 9133 2748
rect 9069 2688 9133 2692
rect 11980 2748 12044 2752
rect 11980 2692 11984 2748
rect 11984 2692 12040 2748
rect 12040 2692 12044 2748
rect 11980 2688 12044 2692
rect 12060 2748 12124 2752
rect 12060 2692 12064 2748
rect 12064 2692 12120 2748
rect 12120 2692 12124 2748
rect 12060 2688 12124 2692
rect 12140 2748 12204 2752
rect 12140 2692 12144 2748
rect 12144 2692 12200 2748
rect 12200 2692 12204 2748
rect 12140 2688 12204 2692
rect 12220 2748 12284 2752
rect 12220 2692 12224 2748
rect 12224 2692 12280 2748
rect 12280 2692 12284 2748
rect 12220 2688 12284 2692
rect 3187 2204 3251 2208
rect 3187 2148 3191 2204
rect 3191 2148 3247 2204
rect 3247 2148 3251 2204
rect 3187 2144 3251 2148
rect 3267 2204 3331 2208
rect 3267 2148 3271 2204
rect 3271 2148 3327 2204
rect 3327 2148 3331 2204
rect 3267 2144 3331 2148
rect 3347 2204 3411 2208
rect 3347 2148 3351 2204
rect 3351 2148 3407 2204
rect 3407 2148 3411 2204
rect 3347 2144 3411 2148
rect 3427 2204 3491 2208
rect 3427 2148 3431 2204
rect 3431 2148 3487 2204
rect 3487 2148 3491 2204
rect 3427 2144 3491 2148
rect 6338 2204 6402 2208
rect 6338 2148 6342 2204
rect 6342 2148 6398 2204
rect 6398 2148 6402 2204
rect 6338 2144 6402 2148
rect 6418 2204 6482 2208
rect 6418 2148 6422 2204
rect 6422 2148 6478 2204
rect 6478 2148 6482 2204
rect 6418 2144 6482 2148
rect 6498 2204 6562 2208
rect 6498 2148 6502 2204
rect 6502 2148 6558 2204
rect 6558 2148 6562 2204
rect 6498 2144 6562 2148
rect 6578 2204 6642 2208
rect 6578 2148 6582 2204
rect 6582 2148 6638 2204
rect 6638 2148 6642 2204
rect 6578 2144 6642 2148
rect 9489 2204 9553 2208
rect 9489 2148 9493 2204
rect 9493 2148 9549 2204
rect 9549 2148 9553 2204
rect 9489 2144 9553 2148
rect 9569 2204 9633 2208
rect 9569 2148 9573 2204
rect 9573 2148 9629 2204
rect 9629 2148 9633 2204
rect 9569 2144 9633 2148
rect 9649 2204 9713 2208
rect 9649 2148 9653 2204
rect 9653 2148 9709 2204
rect 9709 2148 9713 2204
rect 9649 2144 9713 2148
rect 9729 2204 9793 2208
rect 9729 2148 9733 2204
rect 9733 2148 9789 2204
rect 9789 2148 9793 2204
rect 9729 2144 9793 2148
rect 12640 2204 12704 2208
rect 12640 2148 12644 2204
rect 12644 2148 12700 2204
rect 12700 2148 12704 2204
rect 12640 2144 12704 2148
rect 12720 2204 12784 2208
rect 12720 2148 12724 2204
rect 12724 2148 12780 2204
rect 12780 2148 12784 2204
rect 12720 2144 12784 2148
rect 12800 2204 12864 2208
rect 12800 2148 12804 2204
rect 12804 2148 12860 2204
rect 12860 2148 12864 2204
rect 12800 2144 12864 2148
rect 12880 2204 12944 2208
rect 12880 2148 12884 2204
rect 12884 2148 12940 2204
rect 12940 2148 12944 2204
rect 12880 2144 12944 2148
<< metal4 >>
rect 2519 14720 2839 14736
rect 2519 14656 2527 14720
rect 2591 14656 2607 14720
rect 2671 14656 2687 14720
rect 2751 14656 2767 14720
rect 2831 14656 2839 14720
rect 2519 13632 2839 14656
rect 2519 13568 2527 13632
rect 2591 13568 2607 13632
rect 2671 13568 2687 13632
rect 2751 13568 2767 13632
rect 2831 13568 2839 13632
rect 2519 13238 2839 13568
rect 2519 13002 2561 13238
rect 2797 13002 2839 13238
rect 2519 12544 2839 13002
rect 2519 12480 2527 12544
rect 2591 12480 2607 12544
rect 2671 12480 2687 12544
rect 2751 12480 2767 12544
rect 2831 12480 2839 12544
rect 2519 11456 2839 12480
rect 2519 11392 2527 11456
rect 2591 11392 2607 11456
rect 2671 11392 2687 11456
rect 2751 11392 2767 11456
rect 2831 11392 2839 11456
rect 2519 10368 2839 11392
rect 2519 10304 2527 10368
rect 2591 10304 2607 10368
rect 2671 10304 2687 10368
rect 2751 10304 2767 10368
rect 2831 10304 2839 10368
rect 2519 10111 2839 10304
rect 2519 9875 2561 10111
rect 2797 9875 2839 10111
rect 2519 9280 2839 9875
rect 2519 9216 2527 9280
rect 2591 9216 2607 9280
rect 2671 9216 2687 9280
rect 2751 9216 2767 9280
rect 2831 9216 2839 9280
rect 2519 8192 2839 9216
rect 2519 8128 2527 8192
rect 2591 8128 2607 8192
rect 2671 8128 2687 8192
rect 2751 8128 2767 8192
rect 2831 8128 2839 8192
rect 2519 7104 2839 8128
rect 2519 7040 2527 7104
rect 2591 7040 2607 7104
rect 2671 7040 2687 7104
rect 2751 7040 2767 7104
rect 2831 7040 2839 7104
rect 2519 6984 2839 7040
rect 2519 6748 2561 6984
rect 2797 6748 2839 6984
rect 2519 6016 2839 6748
rect 2519 5952 2527 6016
rect 2591 5952 2607 6016
rect 2671 5952 2687 6016
rect 2751 5952 2767 6016
rect 2831 5952 2839 6016
rect 2519 4928 2839 5952
rect 2519 4864 2527 4928
rect 2591 4864 2607 4928
rect 2671 4864 2687 4928
rect 2751 4864 2767 4928
rect 2831 4864 2839 4928
rect 2519 3857 2839 4864
rect 2519 3840 2561 3857
rect 2797 3840 2839 3857
rect 2519 3776 2527 3840
rect 2831 3776 2839 3840
rect 2519 3621 2561 3776
rect 2797 3621 2839 3776
rect 2519 2752 2839 3621
rect 2519 2688 2527 2752
rect 2591 2688 2607 2752
rect 2671 2688 2687 2752
rect 2751 2688 2767 2752
rect 2831 2688 2839 2752
rect 2519 2128 2839 2688
rect 3179 14176 3499 14736
rect 3179 14112 3187 14176
rect 3251 14112 3267 14176
rect 3331 14112 3347 14176
rect 3411 14112 3427 14176
rect 3491 14112 3499 14176
rect 3179 13898 3499 14112
rect 3179 13662 3221 13898
rect 3457 13662 3499 13898
rect 3179 13088 3499 13662
rect 3179 13024 3187 13088
rect 3251 13024 3267 13088
rect 3331 13024 3347 13088
rect 3411 13024 3427 13088
rect 3491 13024 3499 13088
rect 3179 12000 3499 13024
rect 3179 11936 3187 12000
rect 3251 11936 3267 12000
rect 3331 11936 3347 12000
rect 3411 11936 3427 12000
rect 3491 11936 3499 12000
rect 3179 10912 3499 11936
rect 3179 10848 3187 10912
rect 3251 10848 3267 10912
rect 3331 10848 3347 10912
rect 3411 10848 3427 10912
rect 3491 10848 3499 10912
rect 3179 10771 3499 10848
rect 3179 10535 3221 10771
rect 3457 10535 3499 10771
rect 3179 9824 3499 10535
rect 3179 9760 3187 9824
rect 3251 9760 3267 9824
rect 3331 9760 3347 9824
rect 3411 9760 3427 9824
rect 3491 9760 3499 9824
rect 3179 8736 3499 9760
rect 3179 8672 3187 8736
rect 3251 8672 3267 8736
rect 3331 8672 3347 8736
rect 3411 8672 3427 8736
rect 3491 8672 3499 8736
rect 3179 7648 3499 8672
rect 3179 7584 3187 7648
rect 3251 7644 3267 7648
rect 3331 7644 3347 7648
rect 3411 7644 3427 7648
rect 3491 7584 3499 7648
rect 3179 7408 3221 7584
rect 3457 7408 3499 7584
rect 3179 6560 3499 7408
rect 3179 6496 3187 6560
rect 3251 6496 3267 6560
rect 3331 6496 3347 6560
rect 3411 6496 3427 6560
rect 3491 6496 3499 6560
rect 3179 5472 3499 6496
rect 3179 5408 3187 5472
rect 3251 5408 3267 5472
rect 3331 5408 3347 5472
rect 3411 5408 3427 5472
rect 3491 5408 3499 5472
rect 3179 4517 3499 5408
rect 3179 4384 3221 4517
rect 3457 4384 3499 4517
rect 3179 4320 3187 4384
rect 3491 4320 3499 4384
rect 3179 4281 3221 4320
rect 3457 4281 3499 4320
rect 3179 3296 3499 4281
rect 3179 3232 3187 3296
rect 3251 3232 3267 3296
rect 3331 3232 3347 3296
rect 3411 3232 3427 3296
rect 3491 3232 3499 3296
rect 3179 2208 3499 3232
rect 3179 2144 3187 2208
rect 3251 2144 3267 2208
rect 3331 2144 3347 2208
rect 3411 2144 3427 2208
rect 3491 2144 3499 2208
rect 3179 2128 3499 2144
rect 5670 14720 5990 14736
rect 5670 14656 5678 14720
rect 5742 14656 5758 14720
rect 5822 14656 5838 14720
rect 5902 14656 5918 14720
rect 5982 14656 5990 14720
rect 5670 13632 5990 14656
rect 5670 13568 5678 13632
rect 5742 13568 5758 13632
rect 5822 13568 5838 13632
rect 5902 13568 5918 13632
rect 5982 13568 5990 13632
rect 5670 13238 5990 13568
rect 5670 13002 5712 13238
rect 5948 13002 5990 13238
rect 5670 12544 5990 13002
rect 5670 12480 5678 12544
rect 5742 12480 5758 12544
rect 5822 12480 5838 12544
rect 5902 12480 5918 12544
rect 5982 12480 5990 12544
rect 5670 11456 5990 12480
rect 6330 14176 6650 14736
rect 6330 14112 6338 14176
rect 6402 14112 6418 14176
rect 6482 14112 6498 14176
rect 6562 14112 6578 14176
rect 6642 14112 6650 14176
rect 6330 13898 6650 14112
rect 6330 13662 6372 13898
rect 6608 13662 6650 13898
rect 6330 13088 6650 13662
rect 6330 13024 6338 13088
rect 6402 13024 6418 13088
rect 6482 13024 6498 13088
rect 6562 13024 6578 13088
rect 6642 13024 6650 13088
rect 6131 12340 6197 12341
rect 6131 12276 6132 12340
rect 6196 12276 6197 12340
rect 6131 12275 6197 12276
rect 5670 11392 5678 11456
rect 5742 11392 5758 11456
rect 5822 11392 5838 11456
rect 5902 11392 5918 11456
rect 5982 11392 5990 11456
rect 5670 10368 5990 11392
rect 5670 10304 5678 10368
rect 5742 10304 5758 10368
rect 5822 10304 5838 10368
rect 5902 10304 5918 10368
rect 5982 10304 5990 10368
rect 5670 10111 5990 10304
rect 5670 9875 5712 10111
rect 5948 9875 5990 10111
rect 5670 9280 5990 9875
rect 6134 9621 6194 12275
rect 6330 12000 6650 13024
rect 6330 11936 6338 12000
rect 6402 11936 6418 12000
rect 6482 11936 6498 12000
rect 6562 11936 6578 12000
rect 6642 11936 6650 12000
rect 6330 10912 6650 11936
rect 6330 10848 6338 10912
rect 6402 10848 6418 10912
rect 6482 10848 6498 10912
rect 6562 10848 6578 10912
rect 6642 10848 6650 10912
rect 6330 10771 6650 10848
rect 6330 10535 6372 10771
rect 6608 10535 6650 10771
rect 6330 9824 6650 10535
rect 6330 9760 6338 9824
rect 6402 9760 6418 9824
rect 6482 9760 6498 9824
rect 6562 9760 6578 9824
rect 6642 9760 6650 9824
rect 6131 9620 6197 9621
rect 6131 9556 6132 9620
rect 6196 9556 6197 9620
rect 6131 9555 6197 9556
rect 5670 9216 5678 9280
rect 5742 9216 5758 9280
rect 5822 9216 5838 9280
rect 5902 9216 5918 9280
rect 5982 9216 5990 9280
rect 5670 8192 5990 9216
rect 5670 8128 5678 8192
rect 5742 8128 5758 8192
rect 5822 8128 5838 8192
rect 5902 8128 5918 8192
rect 5982 8128 5990 8192
rect 5670 7104 5990 8128
rect 5670 7040 5678 7104
rect 5742 7040 5758 7104
rect 5822 7040 5838 7104
rect 5902 7040 5918 7104
rect 5982 7040 5990 7104
rect 5670 6984 5990 7040
rect 5670 6748 5712 6984
rect 5948 6748 5990 6984
rect 5670 6016 5990 6748
rect 5670 5952 5678 6016
rect 5742 5952 5758 6016
rect 5822 5952 5838 6016
rect 5902 5952 5918 6016
rect 5982 5952 5990 6016
rect 5670 4928 5990 5952
rect 5670 4864 5678 4928
rect 5742 4864 5758 4928
rect 5822 4864 5838 4928
rect 5902 4864 5918 4928
rect 5982 4864 5990 4928
rect 5670 3857 5990 4864
rect 5670 3840 5712 3857
rect 5948 3840 5990 3857
rect 5670 3776 5678 3840
rect 5982 3776 5990 3840
rect 5670 3621 5712 3776
rect 5948 3621 5990 3776
rect 5670 2752 5990 3621
rect 5670 2688 5678 2752
rect 5742 2688 5758 2752
rect 5822 2688 5838 2752
rect 5902 2688 5918 2752
rect 5982 2688 5990 2752
rect 5670 2128 5990 2688
rect 6330 8736 6650 9760
rect 6330 8672 6338 8736
rect 6402 8672 6418 8736
rect 6482 8672 6498 8736
rect 6562 8672 6578 8736
rect 6642 8672 6650 8736
rect 6330 7648 6650 8672
rect 6330 7584 6338 7648
rect 6402 7644 6418 7648
rect 6482 7644 6498 7648
rect 6562 7644 6578 7648
rect 6642 7584 6650 7648
rect 6330 7408 6372 7584
rect 6608 7408 6650 7584
rect 6330 6560 6650 7408
rect 6330 6496 6338 6560
rect 6402 6496 6418 6560
rect 6482 6496 6498 6560
rect 6562 6496 6578 6560
rect 6642 6496 6650 6560
rect 6330 5472 6650 6496
rect 6330 5408 6338 5472
rect 6402 5408 6418 5472
rect 6482 5408 6498 5472
rect 6562 5408 6578 5472
rect 6642 5408 6650 5472
rect 6330 4517 6650 5408
rect 6330 4384 6372 4517
rect 6608 4384 6650 4517
rect 6330 4320 6338 4384
rect 6642 4320 6650 4384
rect 6330 4281 6372 4320
rect 6608 4281 6650 4320
rect 6330 3296 6650 4281
rect 6330 3232 6338 3296
rect 6402 3232 6418 3296
rect 6482 3232 6498 3296
rect 6562 3232 6578 3296
rect 6642 3232 6650 3296
rect 6330 2208 6650 3232
rect 6330 2144 6338 2208
rect 6402 2144 6418 2208
rect 6482 2144 6498 2208
rect 6562 2144 6578 2208
rect 6642 2144 6650 2208
rect 6330 2128 6650 2144
rect 8821 14720 9141 14736
rect 8821 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9069 14720
rect 9133 14656 9141 14720
rect 8821 13632 9141 14656
rect 8821 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9069 13632
rect 9133 13568 9141 13632
rect 8821 13238 9141 13568
rect 8821 13002 8863 13238
rect 9099 13002 9141 13238
rect 8821 12544 9141 13002
rect 8821 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9069 12544
rect 9133 12480 9141 12544
rect 8821 11456 9141 12480
rect 8821 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9069 11456
rect 9133 11392 9141 11456
rect 8821 10368 9141 11392
rect 8821 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9069 10368
rect 9133 10304 9141 10368
rect 8821 10111 9141 10304
rect 8821 9875 8863 10111
rect 9099 9875 9141 10111
rect 8821 9280 9141 9875
rect 8821 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9069 9280
rect 9133 9216 9141 9280
rect 8821 8192 9141 9216
rect 8821 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9069 8192
rect 9133 8128 9141 8192
rect 8821 7104 9141 8128
rect 8821 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9069 7104
rect 9133 7040 9141 7104
rect 8821 6984 9141 7040
rect 8821 6748 8863 6984
rect 9099 6748 9141 6984
rect 8821 6016 9141 6748
rect 8821 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9069 6016
rect 9133 5952 9141 6016
rect 8821 4928 9141 5952
rect 8821 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9069 4928
rect 9133 4864 9141 4928
rect 8821 3857 9141 4864
rect 8821 3840 8863 3857
rect 9099 3840 9141 3857
rect 8821 3776 8829 3840
rect 9133 3776 9141 3840
rect 8821 3621 8863 3776
rect 9099 3621 9141 3776
rect 8821 2752 9141 3621
rect 8821 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9069 2752
rect 9133 2688 9141 2752
rect 8821 2128 9141 2688
rect 9481 14176 9801 14736
rect 9481 14112 9489 14176
rect 9553 14112 9569 14176
rect 9633 14112 9649 14176
rect 9713 14112 9729 14176
rect 9793 14112 9801 14176
rect 9481 13898 9801 14112
rect 9481 13662 9523 13898
rect 9759 13662 9801 13898
rect 9481 13088 9801 13662
rect 9481 13024 9489 13088
rect 9553 13024 9569 13088
rect 9633 13024 9649 13088
rect 9713 13024 9729 13088
rect 9793 13024 9801 13088
rect 9481 12000 9801 13024
rect 9481 11936 9489 12000
rect 9553 11936 9569 12000
rect 9633 11936 9649 12000
rect 9713 11936 9729 12000
rect 9793 11936 9801 12000
rect 9481 10912 9801 11936
rect 9481 10848 9489 10912
rect 9553 10848 9569 10912
rect 9633 10848 9649 10912
rect 9713 10848 9729 10912
rect 9793 10848 9801 10912
rect 9481 10771 9801 10848
rect 9481 10535 9523 10771
rect 9759 10535 9801 10771
rect 9481 9824 9801 10535
rect 9481 9760 9489 9824
rect 9553 9760 9569 9824
rect 9633 9760 9649 9824
rect 9713 9760 9729 9824
rect 9793 9760 9801 9824
rect 9481 8736 9801 9760
rect 9481 8672 9489 8736
rect 9553 8672 9569 8736
rect 9633 8672 9649 8736
rect 9713 8672 9729 8736
rect 9793 8672 9801 8736
rect 9481 7648 9801 8672
rect 9481 7584 9489 7648
rect 9553 7644 9569 7648
rect 9633 7644 9649 7648
rect 9713 7644 9729 7648
rect 9793 7584 9801 7648
rect 9481 7408 9523 7584
rect 9759 7408 9801 7584
rect 9481 6560 9801 7408
rect 9481 6496 9489 6560
rect 9553 6496 9569 6560
rect 9633 6496 9649 6560
rect 9713 6496 9729 6560
rect 9793 6496 9801 6560
rect 9481 5472 9801 6496
rect 9481 5408 9489 5472
rect 9553 5408 9569 5472
rect 9633 5408 9649 5472
rect 9713 5408 9729 5472
rect 9793 5408 9801 5472
rect 9481 4517 9801 5408
rect 9481 4384 9523 4517
rect 9759 4384 9801 4517
rect 9481 4320 9489 4384
rect 9793 4320 9801 4384
rect 9481 4281 9523 4320
rect 9759 4281 9801 4320
rect 9481 3296 9801 4281
rect 9481 3232 9489 3296
rect 9553 3232 9569 3296
rect 9633 3232 9649 3296
rect 9713 3232 9729 3296
rect 9793 3232 9801 3296
rect 9481 2208 9801 3232
rect 9481 2144 9489 2208
rect 9553 2144 9569 2208
rect 9633 2144 9649 2208
rect 9713 2144 9729 2208
rect 9793 2144 9801 2208
rect 9481 2128 9801 2144
rect 11972 14720 12292 14736
rect 11972 14656 11980 14720
rect 12044 14656 12060 14720
rect 12124 14656 12140 14720
rect 12204 14656 12220 14720
rect 12284 14656 12292 14720
rect 11972 13632 12292 14656
rect 11972 13568 11980 13632
rect 12044 13568 12060 13632
rect 12124 13568 12140 13632
rect 12204 13568 12220 13632
rect 12284 13568 12292 13632
rect 11972 13238 12292 13568
rect 11972 13002 12014 13238
rect 12250 13002 12292 13238
rect 11972 12544 12292 13002
rect 11972 12480 11980 12544
rect 12044 12480 12060 12544
rect 12124 12480 12140 12544
rect 12204 12480 12220 12544
rect 12284 12480 12292 12544
rect 11972 11456 12292 12480
rect 11972 11392 11980 11456
rect 12044 11392 12060 11456
rect 12124 11392 12140 11456
rect 12204 11392 12220 11456
rect 12284 11392 12292 11456
rect 11972 10368 12292 11392
rect 11972 10304 11980 10368
rect 12044 10304 12060 10368
rect 12124 10304 12140 10368
rect 12204 10304 12220 10368
rect 12284 10304 12292 10368
rect 11972 10111 12292 10304
rect 11972 9875 12014 10111
rect 12250 9875 12292 10111
rect 11972 9280 12292 9875
rect 11972 9216 11980 9280
rect 12044 9216 12060 9280
rect 12124 9216 12140 9280
rect 12204 9216 12220 9280
rect 12284 9216 12292 9280
rect 11972 8192 12292 9216
rect 11972 8128 11980 8192
rect 12044 8128 12060 8192
rect 12124 8128 12140 8192
rect 12204 8128 12220 8192
rect 12284 8128 12292 8192
rect 11972 7104 12292 8128
rect 11972 7040 11980 7104
rect 12044 7040 12060 7104
rect 12124 7040 12140 7104
rect 12204 7040 12220 7104
rect 12284 7040 12292 7104
rect 11972 6984 12292 7040
rect 11972 6748 12014 6984
rect 12250 6748 12292 6984
rect 11972 6016 12292 6748
rect 11972 5952 11980 6016
rect 12044 5952 12060 6016
rect 12124 5952 12140 6016
rect 12204 5952 12220 6016
rect 12284 5952 12292 6016
rect 11972 4928 12292 5952
rect 11972 4864 11980 4928
rect 12044 4864 12060 4928
rect 12124 4864 12140 4928
rect 12204 4864 12220 4928
rect 12284 4864 12292 4928
rect 11972 3857 12292 4864
rect 11972 3840 12014 3857
rect 12250 3840 12292 3857
rect 11972 3776 11980 3840
rect 12284 3776 12292 3840
rect 11972 3621 12014 3776
rect 12250 3621 12292 3776
rect 11972 2752 12292 3621
rect 11972 2688 11980 2752
rect 12044 2688 12060 2752
rect 12124 2688 12140 2752
rect 12204 2688 12220 2752
rect 12284 2688 12292 2752
rect 11972 2128 12292 2688
rect 12632 14176 12952 14736
rect 12632 14112 12640 14176
rect 12704 14112 12720 14176
rect 12784 14112 12800 14176
rect 12864 14112 12880 14176
rect 12944 14112 12952 14176
rect 12632 13898 12952 14112
rect 12632 13662 12674 13898
rect 12910 13662 12952 13898
rect 12632 13088 12952 13662
rect 12632 13024 12640 13088
rect 12704 13024 12720 13088
rect 12784 13024 12800 13088
rect 12864 13024 12880 13088
rect 12944 13024 12952 13088
rect 12632 12000 12952 13024
rect 12632 11936 12640 12000
rect 12704 11936 12720 12000
rect 12784 11936 12800 12000
rect 12864 11936 12880 12000
rect 12944 11936 12952 12000
rect 12632 10912 12952 11936
rect 12632 10848 12640 10912
rect 12704 10848 12720 10912
rect 12784 10848 12800 10912
rect 12864 10848 12880 10912
rect 12944 10848 12952 10912
rect 12632 10771 12952 10848
rect 12632 10535 12674 10771
rect 12910 10535 12952 10771
rect 12632 9824 12952 10535
rect 12632 9760 12640 9824
rect 12704 9760 12720 9824
rect 12784 9760 12800 9824
rect 12864 9760 12880 9824
rect 12944 9760 12952 9824
rect 12632 8736 12952 9760
rect 12632 8672 12640 8736
rect 12704 8672 12720 8736
rect 12784 8672 12800 8736
rect 12864 8672 12880 8736
rect 12944 8672 12952 8736
rect 12632 7648 12952 8672
rect 12632 7584 12640 7648
rect 12704 7644 12720 7648
rect 12784 7644 12800 7648
rect 12864 7644 12880 7648
rect 12944 7584 12952 7648
rect 12632 7408 12674 7584
rect 12910 7408 12952 7584
rect 12632 6560 12952 7408
rect 12632 6496 12640 6560
rect 12704 6496 12720 6560
rect 12784 6496 12800 6560
rect 12864 6496 12880 6560
rect 12944 6496 12952 6560
rect 12632 5472 12952 6496
rect 12632 5408 12640 5472
rect 12704 5408 12720 5472
rect 12784 5408 12800 5472
rect 12864 5408 12880 5472
rect 12944 5408 12952 5472
rect 12632 4517 12952 5408
rect 12632 4384 12674 4517
rect 12910 4384 12952 4517
rect 12632 4320 12640 4384
rect 12944 4320 12952 4384
rect 12632 4281 12674 4320
rect 12910 4281 12952 4320
rect 12632 3296 12952 4281
rect 12632 3232 12640 3296
rect 12704 3232 12720 3296
rect 12784 3232 12800 3296
rect 12864 3232 12880 3296
rect 12944 3232 12952 3296
rect 12632 2208 12952 3232
rect 12632 2144 12640 2208
rect 12704 2144 12720 2208
rect 12784 2144 12800 2208
rect 12864 2144 12880 2208
rect 12944 2144 12952 2208
rect 12632 2128 12952 2144
<< via4 >>
rect 2561 13002 2797 13238
rect 2561 9875 2797 10111
rect 2561 6748 2797 6984
rect 2561 3840 2797 3857
rect 2561 3776 2591 3840
rect 2591 3776 2607 3840
rect 2607 3776 2671 3840
rect 2671 3776 2687 3840
rect 2687 3776 2751 3840
rect 2751 3776 2767 3840
rect 2767 3776 2797 3840
rect 2561 3621 2797 3776
rect 3221 13662 3457 13898
rect 3221 10535 3457 10771
rect 3221 7584 3251 7644
rect 3251 7584 3267 7644
rect 3267 7584 3331 7644
rect 3331 7584 3347 7644
rect 3347 7584 3411 7644
rect 3411 7584 3427 7644
rect 3427 7584 3457 7644
rect 3221 7408 3457 7584
rect 3221 4384 3457 4517
rect 3221 4320 3251 4384
rect 3251 4320 3267 4384
rect 3267 4320 3331 4384
rect 3331 4320 3347 4384
rect 3347 4320 3411 4384
rect 3411 4320 3427 4384
rect 3427 4320 3457 4384
rect 3221 4281 3457 4320
rect 5712 13002 5948 13238
rect 6372 13662 6608 13898
rect 5712 9875 5948 10111
rect 6372 10535 6608 10771
rect 5712 6748 5948 6984
rect 5712 3840 5948 3857
rect 5712 3776 5742 3840
rect 5742 3776 5758 3840
rect 5758 3776 5822 3840
rect 5822 3776 5838 3840
rect 5838 3776 5902 3840
rect 5902 3776 5918 3840
rect 5918 3776 5948 3840
rect 5712 3621 5948 3776
rect 6372 7584 6402 7644
rect 6402 7584 6418 7644
rect 6418 7584 6482 7644
rect 6482 7584 6498 7644
rect 6498 7584 6562 7644
rect 6562 7584 6578 7644
rect 6578 7584 6608 7644
rect 6372 7408 6608 7584
rect 6372 4384 6608 4517
rect 6372 4320 6402 4384
rect 6402 4320 6418 4384
rect 6418 4320 6482 4384
rect 6482 4320 6498 4384
rect 6498 4320 6562 4384
rect 6562 4320 6578 4384
rect 6578 4320 6608 4384
rect 6372 4281 6608 4320
rect 8863 13002 9099 13238
rect 8863 9875 9099 10111
rect 8863 6748 9099 6984
rect 8863 3840 9099 3857
rect 8863 3776 8893 3840
rect 8893 3776 8909 3840
rect 8909 3776 8973 3840
rect 8973 3776 8989 3840
rect 8989 3776 9053 3840
rect 9053 3776 9069 3840
rect 9069 3776 9099 3840
rect 8863 3621 9099 3776
rect 9523 13662 9759 13898
rect 9523 10535 9759 10771
rect 9523 7584 9553 7644
rect 9553 7584 9569 7644
rect 9569 7584 9633 7644
rect 9633 7584 9649 7644
rect 9649 7584 9713 7644
rect 9713 7584 9729 7644
rect 9729 7584 9759 7644
rect 9523 7408 9759 7584
rect 9523 4384 9759 4517
rect 9523 4320 9553 4384
rect 9553 4320 9569 4384
rect 9569 4320 9633 4384
rect 9633 4320 9649 4384
rect 9649 4320 9713 4384
rect 9713 4320 9729 4384
rect 9729 4320 9759 4384
rect 9523 4281 9759 4320
rect 12014 13002 12250 13238
rect 12014 9875 12250 10111
rect 12014 6748 12250 6984
rect 12014 3840 12250 3857
rect 12014 3776 12044 3840
rect 12044 3776 12060 3840
rect 12060 3776 12124 3840
rect 12124 3776 12140 3840
rect 12140 3776 12204 3840
rect 12204 3776 12220 3840
rect 12220 3776 12250 3840
rect 12014 3621 12250 3776
rect 12674 13662 12910 13898
rect 12674 10535 12910 10771
rect 12674 7584 12704 7644
rect 12704 7584 12720 7644
rect 12720 7584 12784 7644
rect 12784 7584 12800 7644
rect 12800 7584 12864 7644
rect 12864 7584 12880 7644
rect 12880 7584 12910 7644
rect 12674 7408 12910 7584
rect 12674 4384 12910 4517
rect 12674 4320 12704 4384
rect 12704 4320 12720 4384
rect 12720 4320 12784 4384
rect 12784 4320 12800 4384
rect 12800 4320 12864 4384
rect 12864 4320 12880 4384
rect 12880 4320 12910 4384
rect 12674 4281 12910 4320
<< metal5 >>
rect 1056 13898 13756 13940
rect 1056 13662 3221 13898
rect 3457 13662 6372 13898
rect 6608 13662 9523 13898
rect 9759 13662 12674 13898
rect 12910 13662 13756 13898
rect 1056 13620 13756 13662
rect 1056 13238 13756 13280
rect 1056 13002 2561 13238
rect 2797 13002 5712 13238
rect 5948 13002 8863 13238
rect 9099 13002 12014 13238
rect 12250 13002 13756 13238
rect 1056 12960 13756 13002
rect 1056 10771 13756 10813
rect 1056 10535 3221 10771
rect 3457 10535 6372 10771
rect 6608 10535 9523 10771
rect 9759 10535 12674 10771
rect 12910 10535 13756 10771
rect 1056 10493 13756 10535
rect 1056 10111 13756 10153
rect 1056 9875 2561 10111
rect 2797 9875 5712 10111
rect 5948 9875 8863 10111
rect 9099 9875 12014 10111
rect 12250 9875 13756 10111
rect 1056 9833 13756 9875
rect 1056 7644 13756 7686
rect 1056 7408 3221 7644
rect 3457 7408 6372 7644
rect 6608 7408 9523 7644
rect 9759 7408 12674 7644
rect 12910 7408 13756 7644
rect 1056 7366 13756 7408
rect 1056 6984 13756 7026
rect 1056 6748 2561 6984
rect 2797 6748 5712 6984
rect 5948 6748 8863 6984
rect 9099 6748 12014 6984
rect 12250 6748 13756 6984
rect 1056 6706 13756 6748
rect 1056 4517 13756 4559
rect 1056 4281 3221 4517
rect 3457 4281 6372 4517
rect 6608 4281 9523 4517
rect 9759 4281 12674 4517
rect 12910 4281 13756 4517
rect 1056 4239 13756 4281
rect 1056 3857 13756 3899
rect 1056 3621 2561 3857
rect 2797 3621 5712 3857
rect 5948 3621 8863 3857
rect 9099 3621 12014 3857
rect 12250 3621 13756 3857
rect 1056 3579 13756 3621
use sky130_fd_sc_hd__and4_2  _175_
timestamp 0
transform -1 0 5704 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _176_
timestamp 0
transform 1 0 3772 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _177_
timestamp 0
transform -1 0 5428 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _178_
timestamp 0
transform -1 0 12788 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_1  _179_
timestamp 0
transform -1 0 9292 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _180_
timestamp 0
transform 1 0 6348 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _181_
timestamp 0
transform -1 0 8096 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _182_
timestamp 0
transform -1 0 11132 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _183_
timestamp 0
transform -1 0 8832 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _184_
timestamp 0
transform 1 0 4784 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _185_
timestamp 0
transform -1 0 7360 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _186_
timestamp 0
transform 1 0 7912 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _187_
timestamp 0
transform 1 0 10580 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _188_
timestamp 0
transform -1 0 12144 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _189_
timestamp 0
transform 1 0 9200 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _190_
timestamp 0
transform -1 0 10580 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_1  _191_
timestamp 0
transform 1 0 8924 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _192_
timestamp 0
transform -1 0 10304 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor3b_1  _193_
timestamp 0
transform -1 0 7084 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nand4_1  _194_
timestamp 0
transform 1 0 8096 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _195_
timestamp 0
transform -1 0 9200 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _196_
timestamp 0
transform 1 0 8188 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _197_
timestamp 0
transform 1 0 8372 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _198_
timestamp 0
transform 1 0 8464 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _199_
timestamp 0
transform -1 0 9200 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _200_
timestamp 0
transform 1 0 10028 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _201_
timestamp 0
transform -1 0 9752 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _202_
timestamp 0
transform -1 0 5888 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _203_
timestamp 0
transform 1 0 8924 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _204_
timestamp 0
transform 1 0 8372 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _205_
timestamp 0
transform -1 0 8924 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _206_
timestamp 0
transform -1 0 10028 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_2  _207_
timestamp 0
transform 1 0 8556 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _208_
timestamp 0
transform 1 0 6440 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _209_
timestamp 0
transform 1 0 5520 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _210_
timestamp 0
transform 1 0 5796 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _211_
timestamp 0
transform -1 0 7084 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _212_
timestamp 0
transform -1 0 6808 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _213_
timestamp 0
transform -1 0 6808 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _214_
timestamp 0
transform -1 0 5888 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _215_
timestamp 0
transform 1 0 5520 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _216_
timestamp 0
transform 1 0 4968 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _217_
timestamp 0
transform -1 0 5060 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _218_
timestamp 0
transform -1 0 3404 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _219_
timestamp 0
transform 1 0 4324 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _220_
timestamp 0
transform 1 0 3680 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _221_
timestamp 0
transform 1 0 4140 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _222_
timestamp 0
transform 1 0 6716 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _223_
timestamp 0
transform -1 0 3772 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _224_
timestamp 0
transform -1 0 3680 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _225_
timestamp 0
transform -1 0 4232 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _226_
timestamp 0
transform -1 0 3036 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _227_
timestamp 0
transform -1 0 1748 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _228_
timestamp 0
transform -1 0 3220 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _229_
timestamp 0
transform 1 0 1840 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _230_
timestamp 0
transform -1 0 2576 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _231_
timestamp 0
transform 1 0 2116 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _232_
timestamp 0
transform 1 0 3772 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _233_
timestamp 0
transform -1 0 3680 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _234_
timestamp 0
transform -1 0 4508 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _235_
timestamp 0
transform -1 0 5152 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _236_
timestamp 0
transform 1 0 4324 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _237_
timestamp 0
transform -1 0 5704 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _238_
timestamp 0
transform 1 0 3864 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _239_
timestamp 0
transform -1 0 3312 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _240_
timestamp 0
transform -1 0 3956 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _241_
timestamp 0
transform -1 0 3036 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _242_
timestamp 0
transform 1 0 2208 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _243_
timestamp 0
transform -1 0 4692 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _244_
timestamp 0
transform -1 0 3588 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _245_
timestamp 0
transform -1 0 3220 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _246_
timestamp 0
transform -1 0 2852 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _247_
timestamp 0
transform 1 0 2116 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _248_
timestamp 0
transform 1 0 3220 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _249_
timestamp 0
transform -1 0 4048 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _250_
timestamp 0
transform -1 0 3312 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _251_
timestamp 0
transform -1 0 2760 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _252_
timestamp 0
transform -1 0 1748 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _253_
timestamp 0
transform 1 0 3772 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _254_
timestamp 0
transform 1 0 4140 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _255_
timestamp 0
transform -1 0 5520 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _256_
timestamp 0
transform -1 0 5060 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _257_
timestamp 0
transform -1 0 4876 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _258_
timestamp 0
transform 1 0 6348 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _259_
timestamp 0
transform -1 0 5980 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _260_
timestamp 0
transform 1 0 4600 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _261_
timestamp 0
transform -1 0 6256 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _262_
timestamp 0
transform -1 0 5152 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _263_
timestamp 0
transform -1 0 4692 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _264_
timestamp 0
transform 1 0 4232 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _265_
timestamp 0
transform -1 0 4232 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _266_
timestamp 0
transform 1 0 3128 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _267_
timestamp 0
transform -1 0 5060 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _268_
timestamp 0
transform 1 0 5520 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _269_
timestamp 0
transform 1 0 4784 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _270_
timestamp 0
transform -1 0 6256 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _271_
timestamp 0
transform 1 0 6348 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _272_
timestamp 0
transform 1 0 6808 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _273_
timestamp 0
transform -1 0 7084 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _274_
timestamp 0
transform 1 0 6072 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _275_
timestamp 0
transform 1 0 6348 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _276_
timestamp 0
transform -1 0 9200 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _277_
timestamp 0
transform -1 0 8556 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _278_
timestamp 0
transform 1 0 7176 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _279_
timestamp 0
transform 1 0 8556 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _280_
timestamp 0
transform 1 0 7636 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _281_
timestamp 0
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _282_
timestamp 0
transform 1 0 7636 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _283_
timestamp 0
transform -1 0 9476 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _284_
timestamp 0
transform 1 0 9292 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _285_
timestamp 0
transform -1 0 9936 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _286_
timestamp 0
transform 1 0 8096 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _287_
timestamp 0
transform -1 0 8832 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _288_
timestamp 0
transform -1 0 8096 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _289_
timestamp 0
transform 1 0 10856 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _290_
timestamp 0
transform 1 0 7360 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _291_
timestamp 0
transform 1 0 8004 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _292_
timestamp 0
transform -1 0 11132 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _293_
timestamp 0
transform 1 0 10120 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_1  _294_
timestamp 0
transform 1 0 11408 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _295_
timestamp 0
transform -1 0 12052 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _296_
timestamp 0
transform 1 0 12052 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _297_
timestamp 0
transform 1 0 12512 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _298_
timestamp 0
transform -1 0 12512 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _299_
timestamp 0
transform -1 0 11868 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _300_
timestamp 0
transform -1 0 12236 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_1  _301_
timestamp 0
transform -1 0 12236 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a41o_1  _302_
timestamp 0
transform 1 0 11408 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _303_
timestamp 0
transform -1 0 11408 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _304_
timestamp 0
transform 1 0 10488 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _305_
timestamp 0
transform 1 0 10948 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _306_
timestamp 0
transform 1 0 11408 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _307_
timestamp 0
transform -1 0 11132 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _308_
timestamp 0
transform 1 0 10488 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _309_
timestamp 0
transform 1 0 9752 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a41o_1  _310_
timestamp 0
transform 1 0 10580 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _311_
timestamp 0
transform -1 0 11408 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _312_
timestamp 0
transform -1 0 10580 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _313_
timestamp 0
transform 1 0 10396 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _314_
timestamp 0
transform -1 0 11408 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _315_
timestamp 0
transform 1 0 9200 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _316_
timestamp 0
transform -1 0 8096 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _317_
timestamp 0
transform 1 0 8188 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _318_
timestamp 0
transform 1 0 7912 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _319_
timestamp 0
transform 1 0 12972 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _320_
timestamp 0
transform -1 0 12696 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _321_
timestamp 0
transform -1 0 7544 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _322_
timestamp 0
transform 1 0 6900 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _323_
timestamp 0
transform 1 0 4048 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _324_
timestamp 0
transform 1 0 3404 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _325_
timestamp 0
transform -1 0 3128 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _326_
timestamp 0
transform -1 0 3404 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _327_
timestamp 0
transform -1 0 6992 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _328_
timestamp 0
transform -1 0 6164 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _329_
timestamp 0
transform -1 0 6624 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _330_
timestamp 0
transform -1 0 2944 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _331_
timestamp 0
transform -1 0 3772 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _332_
timestamp 0
transform -1 0 3036 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _333_
timestamp 0
transform 1 0 7452 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _334_
timestamp 0
transform -1 0 7084 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _335_
timestamp 0
transform 1 0 3404 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _336_
timestamp 0
transform -1 0 7360 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _337_
timestamp 0
transform -1 0 7176 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _338_
timestamp 0
transform 1 0 8004 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _339_
timestamp 0
transform -1 0 10028 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _340_
timestamp 0
transform -1 0 9752 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _341_
timestamp 0
transform -1 0 9752 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _342_
timestamp 0
transform 1 0 10304 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _343_
timestamp 0
transform -1 0 13064 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _344_
timestamp 0
transform 1 0 11960 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _345_
timestamp 0
transform 1 0 12512 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _346_
timestamp 0
transform 1 0 12052 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _347_
timestamp 0
transform -1 0 11408 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _348_
timestamp 0
transform 1 0 13064 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _349_
timestamp 0
transform 1 0 8096 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _350_
timestamp 0
transform -1 0 9844 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _351_
timestamp 0
transform 1 0 8924 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _352_
timestamp 0
transform 1 0 10304 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _353_
timestamp 0
transform 1 0 10764 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _354_
timestamp 0
transform 1 0 5428 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _355_
timestamp 0
transform 1 0 5888 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _356_
timestamp 0
transform 1 0 3128 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _357_
timestamp 0
transform 1 0 3772 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _358_
timestamp 0
transform 1 0 1748 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _359_
timestamp 0
transform 1 0 1472 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _360_
timestamp 0
transform 1 0 4048 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _361_
timestamp 0
transform -1 0 6256 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _362_
timestamp 0
transform 1 0 1656 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _363_
timestamp 0
transform 1 0 1656 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _364_
timestamp 0
transform 1 0 1748 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _365_
timestamp 0
transform 1 0 4876 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _366_
timestamp 0
transform 1 0 5152 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _367_
timestamp 0
transform 1 0 2576 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _368_
timestamp 0
transform 1 0 4416 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _369_
timestamp 0
transform 1 0 5060 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _370_
timestamp 0
transform 1 0 8004 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _371_
timestamp 0
transform -1 0 9844 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _372_
timestamp 0
transform 1 0 7912 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _373_
timestamp 0
transform 1 0 9292 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _374_
timestamp 0
transform 1 0 11500 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _375_
timestamp 0
transform 1 0 11132 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _376_
timestamp 0
transform 1 0 11500 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _377_
timestamp 0
transform 1 0 11500 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _378_
timestamp 0
transform 1 0 9476 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _379_
timestamp 0
transform 1 0 11500 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _380_
timestamp 0
transform 1 0 6992 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 0
transform 1 0 6532 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 0
transform -1 0 6624 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 0
transform 1 0 9108 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 0
transform -1 0 5796 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 0
transform 1 0 8924 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_4  clkload0
timestamp 0
transform 1 0 4784 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  clkload1
timestamp 0
transform 1 0 3956 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  clkload2
timestamp 0
transform 1 0 8924 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3
timestamp 0
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 0
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 0
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_29
timestamp 0
transform 1 0 3772 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_35
timestamp 0
transform 1 0 4324 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_47
timestamp 0
transform 1 0 5428 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_55
timestamp 0
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_57
timestamp 0
transform 1 0 6348 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_65
timestamp 0
transform 1 0 7084 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 0
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 0
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_85
timestamp 0
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_91
timestamp 0
transform 1 0 9476 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_98
timestamp 0
transform 1 0 10120 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_105
timestamp 0
transform 1 0 10764 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_111
timestamp 0
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 0
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_125
timestamp 0
transform 1 0 12604 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_133
timestamp 0
transform 1 0 13340 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_6
timestamp 0
transform 1 0 1656 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_18
timestamp 0
transform 1 0 2760 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_52
timestamp 0
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_62
timestamp 0
transform 1 0 6808 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_66
timestamp 0
transform 1 0 7176 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_74
timestamp 0
transform 1 0 7912 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_100
timestamp 0
transform 1 0 10304 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 0
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_125
timestamp 0
transform 1 0 12604 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_6
timestamp 0
transform 1 0 1656 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_18
timestamp 0
transform 1 0 2760 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_72
timestamp 0
transform 1 0 7728 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_125
timestamp 0
transform 1 0 12604 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 0
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 0
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_27
timestamp 0
transform 1 0 3588 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_50
timestamp 0
transform 1 0 5704 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_54
timestamp 0
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_65
timestamp 0
transform 1 0 7084 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_73
timestamp 0
transform 1 0 7820 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_110
timestamp 0
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_120
timestamp 0
transform 1 0 12144 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_132
timestamp 0
transform 1 0 13248 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 0
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 0
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 0
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_29
timestamp 0
transform 1 0 3772 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_36
timestamp 0
transform 1 0 4416 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_43
timestamp 0
transform 1 0 5060 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_70
timestamp 0
transform 1 0 7544 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_78
timestamp 0
transform 1 0 8280 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_95
timestamp 0
transform 1 0 9844 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_120
timestamp 0
transform 1 0 12144 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_126
timestamp 0
transform 1 0 12696 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_3
timestamp 0
transform 1 0 1380 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_14
timestamp 0
transform 1 0 2392 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_18
timestamp 0
transform 1 0 2760 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_25
timestamp 0
transform 1 0 3404 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_37
timestamp 0
transform 1 0 4508 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_46
timestamp 0
transform 1 0 5336 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_54
timestamp 0
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 0
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 0
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 0
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 0
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 0
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 0
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 0
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_125
timestamp 0
transform 1 0 12604 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_133
timestamp 0
transform 1 0 13340 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_3
timestamp 0
transform 1 0 1380 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_24
timestamp 0
transform 1 0 3312 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_34
timestamp 0
transform 1 0 4232 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_60
timestamp 0
transform 1 0 6624 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_72
timestamp 0
transform 1 0 7728 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_85
timestamp 0
transform 1 0 8924 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_107
timestamp 0
transform 1 0 10948 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_112
timestamp 0
transform 1 0 11408 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_124
timestamp 0
transform 1 0 12512 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_132
timestamp 0
transform 1 0 13248 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_3
timestamp 0
transform 1 0 1380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_27
timestamp 0
transform 1 0 3588 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_44
timestamp 0
transform 1 0 5152 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_57
timestamp 0
transform 1 0 6348 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_62
timestamp 0
transform 1 0 6808 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_79
timestamp 0
transform 1 0 8372 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_100
timestamp 0
transform 1 0 10304 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_3
timestamp 0
transform 1 0 1380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_7
timestamp 0
transform 1 0 1748 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_55
timestamp 0
transform 1 0 6164 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_85
timestamp 0
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_111
timestamp 0
transform 1 0 11316 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 0
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_15
timestamp 0
transform 1 0 2484 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_23
timestamp 0
transform 1 0 3220 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_60
timestamp 0
transform 1 0 6624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_65
timestamp 0
transform 1 0 7084 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_73
timestamp 0
transform 1 0 7820 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_89
timestamp 0
transform 1 0 9292 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 0
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_133
timestamp 0
transform 1 0 13340 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 0
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_15
timestamp 0
transform 1 0 2484 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_20
timestamp 0
transform 1 0 2944 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_29
timestamp 0
transform 1 0 3772 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_50
timestamp 0
transform 1 0 5704 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_62
timestamp 0
transform 1 0 6808 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_85
timestamp 0
transform 1 0 8924 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_116
timestamp 0
transform 1 0 11776 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_128
timestamp 0
transform 1 0 12880 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_3
timestamp 0
transform 1 0 1380 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_31
timestamp 0
transform 1 0 3956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_43
timestamp 0
transform 1 0 5060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 0
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_57
timestamp 0
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_68
timestamp 0
transform 1 0 7360 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_85
timestamp 0
transform 1 0 8924 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_97
timestamp 0
transform 1 0 10028 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_101
timestamp 0
transform 1 0 10396 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 0
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 0
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 0
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_125
timestamp 0
transform 1 0 12604 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_133
timestamp 0
transform 1 0 13340 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_3
timestamp 0
transform 1 0 1380 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_11
timestamp 0
transform 1 0 2116 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_15
timestamp 0
transform 1 0 2484 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_21
timestamp 0
transform 1 0 3036 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 0
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_29
timestamp 0
transform 1 0 3772 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_35
timestamp 0
transform 1 0 4324 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_43
timestamp 0
transform 1 0 5060 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_52
timestamp 0
transform 1 0 5888 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_58
timestamp 0
transform 1 0 6440 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 0
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_97
timestamp 0
transform 1 0 10028 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_109
timestamp 0
transform 1 0 11132 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_122
timestamp 0
transform 1 0 12328 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_133
timestamp 0
transform 1 0 13340 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 0
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_15
timestamp 0
transform 1 0 2484 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_24
timestamp 0
transform 1 0 3312 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_32
timestamp 0
transform 1 0 4048 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_46
timestamp 0
transform 1 0 5336 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_54
timestamp 0
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 0
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_69
timestamp 0
transform 1 0 7452 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_73
timestamp 0
transform 1 0 7820 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_94
timestamp 0
transform 1 0 9752 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_106
timestamp 0
transform 1 0 10856 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_133
timestamp 0
transform 1 0 13340 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_3
timestamp 0
transform 1 0 1380 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_11
timestamp 0
transform 1 0 2116 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_32
timestamp 0
transform 1 0 4048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_72
timestamp 0
transform 1 0 7728 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_94
timestamp 0
transform 1 0 9752 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_106
timestamp 0
transform 1 0 10856 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_127
timestamp 0
transform 1 0 12788 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_133
timestamp 0
transform 1 0 13340 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_3
timestamp 0
transform 1 0 1380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_27
timestamp 0
transform 1 0 3588 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_39
timestamp 0
transform 1 0 4692 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_53
timestamp 0
transform 1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_96
timestamp 0
transform 1 0 9936 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_133
timestamp 0
transform 1 0 13340 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_3
timestamp 0
transform 1 0 1380 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 0
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_29
timestamp 0
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_37
timestamp 0
transform 1 0 4508 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_64
timestamp 0
transform 1 0 6992 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_76
timestamp 0
transform 1 0 8096 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_96
timestamp 0
transform 1 0 9936 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_127
timestamp 0
transform 1 0 12788 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_133
timestamp 0
transform 1 0 13340 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_3
timestamp 0
transform 1 0 1380 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_29
timestamp 0
transform 1 0 3772 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_65
timestamp 0
transform 1 0 7084 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_77
timestamp 0
transform 1 0 8188 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_105
timestamp 0
transform 1 0 10764 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_109
timestamp 0
transform 1 0 11132 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_121
timestamp 0
transform 1 0 12236 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_133
timestamp 0
transform 1 0 13340 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 0
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 0
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 0
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_29
timestamp 0
transform 1 0 3772 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_33
timestamp 0
transform 1 0 4140 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_37
timestamp 0
transform 1 0 4508 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_59
timestamp 0
transform 1 0 6532 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_71
timestamp 0
transform 1 0 7636 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 0
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_85
timestamp 0
transform 1 0 8924 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_129
timestamp 0
transform 1 0 12972 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_133
timestamp 0
transform 1 0 13340 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 0
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_15
timestamp 0
transform 1 0 2484 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_68
timestamp 0
transform 1 0 7360 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_96
timestamp 0
transform 1 0 9936 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_103
timestamp 0
transform 1 0 10580 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 0
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_113
timestamp 0
transform 1 0 11500 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_117
timestamp 0
transform 1 0 11868 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_121
timestamp 0
transform 1 0 12236 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_133
timestamp 0
transform 1 0 13340 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_6
timestamp 0
transform 1 0 1656 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_18
timestamp 0
transform 1 0 2760 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_39
timestamp 0
transform 1 0 4692 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_97
timestamp 0
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_109
timestamp 0
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_121
timestamp 0
transform 1 0 12236 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_129
timestamp 0
transform 1 0 12972 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_6
timestamp 0
transform 1 0 1656 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_18
timestamp 0
transform 1 0 2760 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_30
timestamp 0
transform 1 0 3864 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_42
timestamp 0
transform 1 0 4968 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_48
timestamp 0
transform 1 0 5520 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_60
timestamp 0
transform 1 0 6624 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_72
timestamp 0
transform 1 0 7728 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_95
timestamp 0
transform 1 0 9844 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_107
timestamp 0
transform 1 0 10948 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 0
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_113
timestamp 0
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_125
timestamp 0
transform 1 0 12604 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 0
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 0
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 0
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 0
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_41
timestamp 0
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_53
timestamp 0
transform 1 0 5980 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_57
timestamp 0
transform 1 0 6348 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_69
timestamp 0
transform 1 0 7452 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_81
timestamp 0
transform 1 0 8556 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_85
timestamp 0
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_97
timestamp 0
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_109
timestamp 0
transform 1 0 11132 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_113
timestamp 0
transform 1 0 11500 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_125
timestamp 0
transform 1 0 12604 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_133
timestamp 0
transform 1 0 13340 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 0
transform -1 0 12972 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 0
transform -1 0 10304 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 0
transform -1 0 13340 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 0
transform 1 0 9108 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 0
transform -1 0 7452 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 0
transform 1 0 7176 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output2
timestamp 0
transform -1 0 9476 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output3
timestamp 0
transform -1 0 10120 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output4
timestamp 0
transform -1 0 10764 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output5
timestamp 0
transform 1 0 13064 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_23
timestamp 0
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 0
transform -1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_24
timestamp 0
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 0
transform -1 0 13708 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_25
timestamp 0
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 0
transform -1 0 13708 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_26
timestamp 0
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 0
transform -1 0 13708 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_27
timestamp 0
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 0
transform -1 0 13708 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_28
timestamp 0
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 0
transform -1 0 13708 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_29
timestamp 0
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 0
transform -1 0 13708 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_30
timestamp 0
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 0
transform -1 0 13708 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_31
timestamp 0
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 0
transform -1 0 13708 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_32
timestamp 0
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 0
transform -1 0 13708 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_33
timestamp 0
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 0
transform -1 0 13708 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_34
timestamp 0
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 0
transform -1 0 13708 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_35
timestamp 0
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 0
transform -1 0 13708 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_36
timestamp 0
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 0
transform -1 0 13708 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_37
timestamp 0
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 0
transform -1 0 13708 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_38
timestamp 0
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 0
transform -1 0 13708 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_39
timestamp 0
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 0
transform -1 0 13708 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_40
timestamp 0
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 0
transform -1 0 13708 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_41
timestamp 0
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 0
transform -1 0 13708 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_42
timestamp 0
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 0
transform -1 0 13708 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_43
timestamp 0
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 0
transform -1 0 13708 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_44
timestamp 0
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 0
transform -1 0 13708 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_45
timestamp 0
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 0
transform -1 0 13708 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_46
timestamp 0
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_47
timestamp 0
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_48
timestamp 0
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_49
timestamp 0
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_50
timestamp 0
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_51
timestamp 0
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_52
timestamp 0
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_53
timestamp 0
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_54
timestamp 0
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_55
timestamp 0
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_56
timestamp 0
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_57
timestamp 0
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_58
timestamp 0
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_59
timestamp 0
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_60
timestamp 0
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_61
timestamp 0
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_62
timestamp 0
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_63
timestamp 0
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_64
timestamp 0
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_65
timestamp 0
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_66
timestamp 0
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_67
timestamp 0
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_68
timestamp 0
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_69
timestamp 0
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_70
timestamp 0
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_71
timestamp 0
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_72
timestamp 0
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_73
timestamp 0
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_74
timestamp 0
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_75
timestamp 0
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_76
timestamp 0
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_77
timestamp 0
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_78
timestamp 0
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_79
timestamp 0
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_80
timestamp 0
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_81
timestamp 0
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_82
timestamp 0
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_83
timestamp 0
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_84
timestamp 0
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_85
timestamp 0
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_86
timestamp 0
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_87
timestamp 0
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_88
timestamp 0
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_89
timestamp 0
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_90
timestamp 0
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_91
timestamp 0
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_92
timestamp 0
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_93
timestamp 0
transform 1 0 6256 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_94
timestamp 0
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_95
timestamp 0
transform 1 0 11408 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  ZeroToFiveCounter_6
timestamp 0
transform -1 0 1656 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ZeroToFiveCounter_7
timestamp 0
transform 1 0 13156 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ZeroToFiveCounter_8
timestamp 0
transform -1 0 1656 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ZeroToFiveCounter_9
timestamp 0
transform -1 0 1656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ZeroToFiveCounter_10
timestamp 0
transform 1 0 1380 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ZeroToFiveCounter_11
timestamp 0
transform -1 0 13432 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ZeroToFiveCounter_12
timestamp 0
transform -1 0 13432 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  ZeroToFiveCounter_13
timestamp 0
transform -1 0 13432 0 -1 3264
box -38 -48 314 592
<< labels >>
rlabel metal1 s 7406 14144 7406 14144 4 VGND
rlabel metal1 s 7406 14688 7406 14688 4 VPWR
rlabel metal1 s 5796 4250 5796 4250 4 _000_
rlabel metal1 s 2070 10744 2070 10744 4 _001_
rlabel metal1 s 5014 9962 5014 9962 4 _002_
rlabel metal1 s 5290 11186 5290 11186 4 _003_
rlabel metal2 s 2898 13022 2898 13022 4 _004_
rlabel metal1 s 4784 12410 4784 12410 4 _005_
rlabel metal1 s 5888 13362 5888 13362 4 _006_
rlabel metal1 s 8464 12886 8464 12886 4 _007_
rlabel metal1 s 9476 13498 9476 13498 4 _008_
rlabel metal1 s 8188 9622 8188 9622 4 _009_
rlabel metal1 s 10028 11322 10028 11322 4 _010_
rlabel metal1 s 6026 3434 6026 3434 4 _011_
rlabel metal2 s 12558 7072 12558 7072 4 _012_
rlabel metal1 s 11822 11866 11822 11866 4 _013_
rlabel metal1 s 11592 10574 11592 10574 4 _014_
rlabel metal2 s 11086 9316 11086 9316 4 _015_
rlabel metal1 s 9844 7446 9844 7446 4 _016_
rlabel metal1 s 11592 5882 11592 5882 4 _017_
rlabel metal1 s 9430 6426 9430 6426 4 _018_
rlabel metal1 s 3266 2958 3266 2958 4 _019_
rlabel metal2 s 4140 3434 4140 3434 4 _020_
rlabel metal1 s 1886 6222 1886 6222 4 _021_
rlabel metal1 s 1978 5338 1978 5338 4 _022_
rlabel metal1 s 4416 6426 4416 6426 4 _023_
rlabel metal2 s 5934 7582 5934 7582 4 _024_
rlabel metal2 s 1978 8670 1978 8670 4 _025_
rlabel metal1 s 2070 11322 2070 11322 4 _026_
rlabel metal1 s 8372 3162 8372 3162 4 _027_
rlabel metal1 s 8871 3434 8871 3434 4 _028_
rlabel metal2 s 13110 4284 13110 4284 4 _029_
rlabel metal2 s 12466 3944 12466 3944 4 _030_
rlabel metal1 s 7183 4522 7183 4522 4 _031_
rlabel metal1 s 6992 3162 6992 3162 4 _032_
rlabel metal2 s 4186 2856 4186 2856 4 _033_
rlabel metal1 s 3864 3366 3864 3366 4 _034_
rlabel metal1 s 3036 5338 3036 5338 4 _035_
rlabel metal1 s 3082 5270 3082 5270 4 _036_
rlabel metal1 s 5803 6698 5803 6698 4 _037_
rlabel metal1 s 6118 7514 6118 7514 4 _038_
rlabel metal1 s 2898 8058 2898 8058 4 _039_
rlabel metal1 s 3411 11798 3411 11798 4 _040_
rlabel metal1 s 2990 9622 2990 9622 4 _041_
rlabel metal1 s 6999 9962 6999 9962 4 _042_
rlabel metal1 s 6769 11118 6769 11118 4 _043_
rlabel metal2 s 3542 13022 3542 13022 4 _044_
rlabel metal1 s 6302 12920 6302 12920 4 _045_
rlabel metal1 s 6815 13226 6815 13226 4 _046_
rlabel metal2 s 9890 13022 9890 13022 4 _047_
rlabel metal2 s 9614 13736 9614 13736 4 _048_
rlabel metal1 s 9430 9962 9430 9962 4 _049_
rlabel metal1 s 10396 12614 10396 12614 4 _050_
rlabel metal2 s 12926 6970 12926 6970 4 _051_
rlabel metal1 s 12282 12614 12282 12614 4 _052_
rlabel metal2 s 12558 10846 12558 10846 4 _053_
rlabel metal1 s 12282 9146 12282 9146 4 _054_
rlabel metal2 s 11270 7582 11270 7582 4 _055_
rlabel metal1 s 13117 6358 13117 6358 4 _056_
rlabel metal1 s 8280 6426 8280 6426 4 _057_
rlabel metal1 s 9338 4046 9338 4046 4 _058_
rlabel metal1 s 8960 3706 8960 3706 4 _059_
rlabel metal1 s 10534 4522 10534 4522 4 _060_
rlabel metal1 s 11316 3570 11316 3570 4 _061_
rlabel metal1 s 6808 12614 6808 12614 4 _062_
rlabel metal2 s 7682 8551 7682 8551 4 _063_
rlabel metal1 s 9062 6120 9062 6120 4 _064_
rlabel metal1 s 8464 7786 8464 7786 4 _065_
rlabel metal2 s 5382 9146 5382 9146 4 _066_
rlabel metal1 s 7820 7718 7820 7718 4 _067_
rlabel metal1 s 8418 4624 8418 4624 4 _068_
rlabel metal2 s 11178 3468 11178 3468 4 _069_
rlabel metal2 s 9338 3638 9338 3638 4 _070_
rlabel metal1 s 9384 3162 9384 3162 4 _071_
rlabel metal1 s 9798 3162 9798 3162 4 _072_
rlabel metal1 s 7866 8466 7866 8466 4 _073_
rlabel metal1 s 8602 6222 8602 6222 4 _074_
rlabel metal2 s 8510 4828 8510 4828 4 _075_
rlabel metal2 s 8702 3162 8702 3162 4 _076_
rlabel metal1 s 9062 3162 9062 3162 4 _077_
rlabel metal3 s 9614 6307 9614 6307 4 _078_
rlabel metal2 s 9982 7701 9982 7701 4 _079_
rlabel metal1 s 8510 8466 8510 8466 4 _080_
rlabel metal1 s 8786 10030 8786 10030 4 _081_
rlabel metal1 s 8878 8568 8878 8568 4 _082_
rlabel metal1 s 8878 7310 8878 7310 4 _083_
rlabel metal1 s 9706 6426 9706 6426 4 _084_
rlabel metal1 s 4416 4794 4416 4794 4 _085_
rlabel metal1 s 6670 6392 6670 6392 4 _086_
rlabel metal2 s 6026 4556 6026 4556 4 _087_
rlabel metal1 s 6854 4182 6854 4182 4 _088_
rlabel metal1 s 6302 3162 6302 3162 4 _089_
rlabel metal1 s 5750 3502 5750 3502 4 _090_
rlabel metal1 s 5014 4488 5014 4488 4 _091_
rlabel metal1 s 4968 3162 4968 3162 4 _092_
rlabel metal1 s 3174 3604 3174 3604 4 _093_
rlabel metal1 s 4370 4114 4370 4114 4 _094_
rlabel metal1 s 4324 4250 4324 4250 4 _095_
rlabel metal2 s 2438 10506 2438 10506 4 _096_
rlabel metal2 s 1886 6426 1886 6426 4 _097_
rlabel metal1 s 3266 5746 3266 5746 4 _098_
rlabel metal1 s 3680 5882 3680 5882 4 _099_
rlabel metal1 s 2530 6766 2530 6766 4 _100_
rlabel metal2 s 2346 7072 2346 7072 4 _101_
rlabel metal1 s 2195 6630 2195 6630 4 _102_
rlabel metal1 s 2254 5202 2254 5202 4 _103_
rlabel metal2 s 4186 6460 4186 6460 4 _104_
rlabel metal1 s 3956 6290 3956 6290 4 _105_
rlabel metal1 s 4922 6426 4922 6426 4 _106_
rlabel metal1 s 5474 7888 5474 7888 4 _107_
rlabel metal1 s 3818 9996 3818 9996 4 _108_
rlabel metal1 s 2990 9146 2990 9146 4 _109_
rlabel metal2 s 3542 8704 3542 8704 4 _110_
rlabel metal1 s 2530 8942 2530 8942 4 _111_
rlabel metal1 s 3864 11118 3864 11118 4 _112_
rlabel metal1 s 3036 11322 3036 11322 4 _113_
rlabel metal1 s 2714 11084 2714 11084 4 _114_
rlabel metal1 s 2392 11118 2392 11118 4 _115_
rlabel metal1 s 4002 10064 4002 10064 4 _116_
rlabel metal1 s 2530 10200 2530 10200 4 _117_
rlabel metal2 s 2898 10438 2898 10438 4 _118_
rlabel metal1 s 1932 10234 1932 10234 4 _119_
rlabel metal2 s 4462 10268 4462 10268 4 _120_
rlabel metal2 s 5290 10166 5290 10166 4 _121_
rlabel metal1 s 5336 10778 5336 10778 4 _122_
rlabel metal2 s 4370 10234 4370 10234 4 _123_
rlabel metal1 s 6394 11526 6394 11526 4 _124_
rlabel metal1 s 6118 12206 6118 12206 4 _125_
rlabel metal2 s 5198 11764 5198 11764 4 _126_
rlabel metal2 s 4922 11322 4922 11322 4 _127_
rlabel metal1 s 4140 13498 4140 13498 4 _128_
rlabel metal1 s 4178 13158 4178 13158 4 _129_
rlabel metal1 s 3358 13260 3358 13260 4 _130_
rlabel metal1 s 5014 13158 5014 13158 4 _131_
rlabel metal1 s 5290 12240 5290 12240 4 _132_
rlabel metal1 s 6256 12410 6256 12410 4 _133_
rlabel metal1 s 7038 10506 7038 10506 4 _134_
rlabel metal1 s 7728 12818 7728 12818 4 _135_
rlabel metal1 s 6640 12138 6640 12138 4 _136_
rlabel metal1 s 6670 13906 6670 13906 4 _137_
rlabel metal1 s 8510 13498 8510 13498 4 _138_
rlabel metal1 s 7514 13226 7514 13226 4 _139_
rlabel metal1 s 8786 13328 8786 13328 4 _140_
rlabel metal2 s 7866 13226 7866 13226 4 _141_
rlabel metal1 s 8066 13226 8066 13226 4 _142_
rlabel metal1 s 9246 13362 9246 13362 4 _143_
rlabel metal2 s 8602 9792 8602 9792 4 _144_
rlabel metal1 s 8096 10778 8096 10778 4 _145_
rlabel metal1 s 10718 8908 10718 8908 4 _146_
rlabel metal2 s 8418 9520 8418 9520 4 _147_
rlabel metal2 s 10902 7310 10902 7310 4 _148_
rlabel metal1 s 8004 10642 8004 10642 4 _149_
rlabel metal2 s 8234 10778 8234 10778 4 _150_
rlabel metal1 s 11408 11662 11408 11662 4 _151_
rlabel metal2 s 12282 7446 12282 7446 4 _152_
rlabel metal1 s 12152 7514 12152 7514 4 _153_
rlabel metal1 s 12604 7378 12604 7378 4 _154_
rlabel metal2 s 12374 11526 12374 11526 4 _155_
rlabel metal1 s 11776 11322 11776 11322 4 _156_
rlabel metal1 s 11132 10642 11132 10642 4 _157_
rlabel metal1 s 11362 10234 11362 10234 4 _158_
rlabel metal1 s 10120 7990 10120 7990 4 _159_
rlabel metal1 s 11730 9044 11730 9044 4 _160_
rlabel metal1 s 10626 8976 10626 8976 4 _161_
rlabel metal1 s 10258 7888 10258 7888 4 _162_
rlabel metal2 s 10626 6358 10626 6358 4 _163_
rlabel metal2 s 11270 6698 11270 6698 4 _164_
rlabel metal1 s 10266 6426 10266 6426 4 _165_
rlabel metal1 s 10994 5678 10994 5678 4 _166_
rlabel metal1 s 3864 2414 3864 2414 4 _167_
rlabel metal1 s 3588 13294 3588 13294 4 _168_
rlabel metal1 s 13018 7412 13018 7412 4 _169_
rlabel metal1 s 4048 3978 4048 3978 4 _170_
rlabel metal2 s 5198 7684 5198 7684 4 _171_
rlabel metal1 s 8234 7990 8234 7990 4 _172_
rlabel metal1 s 10534 8500 10534 8500 4 _173_
rlabel metal1 s 8142 10506 8142 10506 4 _174_
rlabel metal4 s 6164 10948 6164 10948 4 clk
rlabel metal1 s 7636 11798 7636 11798 4 clknet_0_clk
rlabel metal1 s 1794 6324 1794 6324 4 clknet_2_0__leaf_clk
rlabel metal2 s 9522 7072 9522 7072 4 clknet_2_1__leaf_clk
rlabel metal1 s 1748 10574 1748 10574 4 clknet_2_2__leaf_clk
rlabel metal1 s 8050 12716 8050 12716 4 clknet_2_3__leaf_clk
rlabel metal2 s 9062 1520 9062 1520 4 count[0]
rlabel metal2 s 9706 959 9706 959 4 count[1]
rlabel metal2 s 10350 1520 10350 1520 4 count[2]
rlabel metal2 s 13294 4301 13294 4301 4 count[3]
rlabel metal1 s 7728 6290 7728 6290 4 net1
rlabel metal3 s 0 12928 800 13048 4 net10
port 2 nsew
rlabel metal2 s 13386 13073 13386 13073 4 net11
rlabel metal2 s 13386 13753 13386 13753 4 net12
rlabel metal2 s 13386 2873 13386 2873 4 net13
rlabel metal1 s 12098 4114 12098 4114 4 net14
rlabel metal1 s 8510 3502 8510 3502 4 net15
rlabel metal1 s 12282 9010 12282 9010 4 net16
rlabel metal2 s 10074 6460 10074 6460 4 net17
rlabel metal1 s 4692 10030 4692 10030 4 net18
rlabel metal1 s 9430 4590 9430 4590 4 net2
rlabel metal1 s 10166 2414 10166 2414 4 net3
rlabel metal1 s 10764 2414 10764 2414 4 net4
rlabel metal1 s 12834 4012 12834 4012 4 net5
rlabel metal3 s 0 2728 800 2848 4 net6
port 1 nsew
rlabel metal3 s 13386 3485 13386 3485 4 net7
rlabel metal3 s 1050 13668 1050 13668 4 net8
rlabel metal3 s 0 3408 800 3528 4 net9
port 6 nsew
rlabel metal2 s 6854 4420 6854 4420 4 one_second_counter\[0\]
rlabel metal1 s 4048 10438 4048 10438 4 one_second_counter\[10\]
rlabel metal2 s 5382 10132 5382 10132 4 one_second_counter\[11\]
rlabel metal2 s 6854 8738 6854 8738 4 one_second_counter\[12\]
rlabel metal1 s 6394 12852 6394 12852 4 one_second_counter\[13\]
rlabel metal1 s 5934 13804 5934 13804 4 one_second_counter\[14\]
rlabel metal1 s 6670 13498 6670 13498 4 one_second_counter\[15\]
rlabel metal1 s 9614 12614 9614 12614 4 one_second_counter\[16\]
rlabel metal2 s 7958 13260 7958 13260 4 one_second_counter\[17\]
rlabel metal1 s 9798 10608 9798 10608 4 one_second_counter\[18\]
rlabel metal2 s 10902 11594 10902 11594 4 one_second_counter\[19\]
rlabel metal1 s 5060 4182 5060 4182 4 one_second_counter\[1\]
rlabel metal2 s 13294 7072 13294 7072 4 one_second_counter\[20\]
rlabel metal1 s 12466 11152 12466 11152 4 one_second_counter\[21\]
rlabel metal1 s 11638 9996 11638 9996 4 one_second_counter\[22\]
rlabel metal2 s 13294 9758 13294 9758 4 one_second_counter\[23\]
rlabel metal1 s 10994 7990 10994 7990 4 one_second_counter\[24\]
rlabel metal1 s 11362 6358 11362 6358 4 one_second_counter\[25\]
rlabel metal2 s 9246 6834 9246 6834 4 one_second_counter\[26\]
rlabel metal1 s 5382 4080 5382 4080 4 one_second_counter\[2\]
rlabel metal2 s 5290 3910 5290 3910 4 one_second_counter\[3\]
rlabel metal1 s 3772 6086 3772 6086 4 one_second_counter\[4\]
rlabel metal2 s 2714 6851 2714 6851 4 one_second_counter\[5\]
rlabel metal1 s 5336 6290 5336 6290 4 one_second_counter\[6\]
rlabel metal1 s 4554 7174 4554 7174 4 one_second_counter\[7\]
rlabel metal1 s 4646 9418 4646 9418 4 one_second_counter\[8\]
rlabel metal1 s 4738 10574 4738 10574 4 one_second_counter\[9\]
rlabel metal2 s 7130 1588 7130 1588 4 rst
flabel metal3 s 400 2788 400 2788 0 FreeSans 600 0 0 0 AN[0]
flabel metal3 s 400 12988 400 12988 0 FreeSans 600 0 0 0 AN[1]
flabel metal3 s 14087 12928 14887 13048 0 FreeSans 600 0 0 0 AN[2]
port 3 nsew
flabel metal3 s 14087 3408 14887 3528 0 FreeSans 600 0 0 0 AN[3]
port 4 nsew
flabel metal3 s 0 13608 800 13728 0 FreeSans 600 0 0 0 AN[4]
port 5 nsew
flabel metal3 s 400 3468 400 3468 0 FreeSans 600 0 0 0 AN[5]
flabel metal3 s 14087 13608 14887 13728 0 FreeSans 600 0 0 0 AN[6]
port 7 nsew
flabel metal3 s 14087 2728 14887 2848 0 FreeSans 600 0 0 0 AN[7]
port 8 nsew
flabel metal5 s 1056 13620 13756 13940 0 FreeSans 3200 0 0 0 VGND
port 9 nsew
flabel metal5 s 1056 10493 13756 10813 0 FreeSans 3200 0 0 0 VGND
port 9 nsew
flabel metal5 s 1056 7366 13756 7686 0 FreeSans 3200 0 0 0 VGND
port 9 nsew
flabel metal5 s 1056 4239 13756 4559 0 FreeSans 3200 0 0 0 VGND
port 9 nsew
flabel metal4 s 12632 2128 12952 14736 0 FreeSans 2400 90 0 0 VGND
port 9 nsew
flabel metal4 s 9481 2128 9801 14736 0 FreeSans 2400 90 0 0 VGND
port 9 nsew
flabel metal4 s 6330 2128 6650 14736 0 FreeSans 2400 90 0 0 VGND
port 9 nsew
flabel metal4 s 3179 2128 3499 14736 0 FreeSans 2400 90 0 0 VGND
port 9 nsew
flabel metal5 s 1056 12960 13756 13280 0 FreeSans 3200 0 0 0 VPWR
port 10 nsew
flabel metal5 s 1056 9833 13756 10153 0 FreeSans 3200 0 0 0 VPWR
port 10 nsew
flabel metal5 s 1056 6706 13756 7026 0 FreeSans 3200 0 0 0 VPWR
port 10 nsew
flabel metal5 s 1056 3579 13756 3899 0 FreeSans 3200 0 0 0 VPWR
port 10 nsew
flabel metal4 s 11972 2128 12292 14736 0 FreeSans 2400 90 0 0 VPWR
port 10 nsew
flabel metal4 s 8821 2128 9141 14736 0 FreeSans 2400 90 0 0 VPWR
port 10 nsew
flabel metal4 s 5670 2128 5990 14736 0 FreeSans 2400 90 0 0 VPWR
port 10 nsew
flabel metal4 s 2519 2128 2839 14736 0 FreeSans 2400 90 0 0 VPWR
port 10 nsew
flabel metal3 s 0 12248 800 12368 0 FreeSans 600 0 0 0 clk
port 11 nsew
flabel metal2 s 9034 0 9090 800 0 FreeSans 280 90 0 0 count[0]
port 12 nsew
flabel metal2 s 9678 0 9734 800 0 FreeSans 280 90 0 0 count[1]
port 13 nsew
flabel metal2 s 10322 0 10378 800 0 FreeSans 280 90 0 0 count[2]
port 14 nsew
flabel metal3 s 14087 4088 14887 4208 0 FreeSans 600 0 0 0 count[3]
port 15 nsew
flabel metal2 s 7102 0 7158 800 0 FreeSans 280 90 0 0 rst
port 16 nsew
<< properties >>
string FIXED_BBOX 0 0 14887 17031
<< end >>
