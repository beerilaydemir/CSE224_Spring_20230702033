* NGSPICE file created from TopModule.ext - technology: sky130A

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

.subckt TopModule Result[13] Result[14] Result[15] Result[16] Result[17] Result[18]
+ Result[19] Result[6] Result[7] Result[8] VGND VPWR clk control reset Result[5] Result[4]
+ Result[3] Result[28] Result[2] Result[27] Result[0] Result[1] Result[26] Result[25]
+ Result[24] Result[12] Result[23] Result[11] Result[22] Result[10] Result[21] Result[9]
+ Result[31] Result[20] Result[30] Result[29]
XFILLER_0_89_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_65_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_484 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_18_Left_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_27_Left_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_36_Left_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_45_Left_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_54_Left_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_63_Left_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_72_Left_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_35_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_81_Left_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_3_Left_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_83_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_59_Right_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_68_Right_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_77_Right_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_86_Right_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_33_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_4_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_78_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_46_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_80_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_51_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_14_Left_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_23_Left_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_32_Left_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_41_Left_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_50_Left_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_7_Left_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_46_Right_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_55_Right_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_64_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_64_Right_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_79_Left_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_73_Right_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_88_Left_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_82_Right_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_16 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_38_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_64_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_75_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTopModule_1 VGND VGND VPWR VPWR TopModule_1/HI Result[0] sky130_fd_sc_hd__conb_1
XFILLER_0_61_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_38_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_10_Left_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_3_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTopModule_2 VGND VGND VPWR VPWR TopModule_2/HI Result[1] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_82_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_54_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_39_Left_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_48_Left_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_42_Right_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_57_Left_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_51_Right_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_66_Left_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_60_Right_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_75_Left_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_84_Left_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_69_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_72_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_89_Right_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTopModule_3 VGND VGND VPWR VPWR TopModule_3/HI Result[2] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_54_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_51_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_67_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_6_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTopModule_4 VGND VGND VPWR VPWR TopModule_4/HI Result[3] sky130_fd_sc_hd__conb_1
XFILLER_0_46_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_2_Left_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_67_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_88_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTopModule_5 VGND VGND VPWR VPWR TopModule_5/HI Result[4] sky130_fd_sc_hd__conb_1
XFILLER_0_34_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_53_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_67_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_17_Left_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_26_Left_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_35_Left_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Left_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_53_Left_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_32_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_62_Left_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_71_Left_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_80_Left_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_74_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_85_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_49_Right_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_58_Right_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTopModule_6 VGND VGND VPWR VPWR TopModule_6/HI Result[5] sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_67_Right_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_76_Right_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_85_Right_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_48_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTopModule_7 VGND VGND VPWR VPWR TopModule_7/HI Result[6] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_3_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Left_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_88_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_71_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTopModule_8 VGND VGND VPWR VPWR TopModule_8/HI Result[7] sky130_fd_sc_hd__conb_1
XFILLER_0_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_67_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_13_Left_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_22_Left_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_32_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_31_Left_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_40_Left_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_88_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_79_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_34_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_6_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_82_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTopModule_9 VGND VGND VPWR VPWR TopModule_9/HI Result[8] sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_45_Right_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_54_Right_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_69_Left_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_63_Right_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_78_Left_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_72_Right_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_87_Left_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_81_Right_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_67_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_88_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_85_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_69_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_79_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_5_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_84_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_2_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_53_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_29_Left_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_38_Left_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_47_Left_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_56_Left_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_50_Right_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_65_Left_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_74_Left_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_83_Left_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_1_Left_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_32_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_79_Right_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_88_Right_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_19_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_16_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_13_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_77_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_79_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_16_Left_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_50_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_25_Left_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_34_Left_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_43_Left_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_52_Left_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_61_Left_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_70_Left_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Left_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_89_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_48_Right_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_57_Right_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_87_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_66_Right_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_75_Right_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_84_Right_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_5_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_47_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_172 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_31_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_73_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_12_Left_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_21_Left_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_30_Left_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_63_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_60_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_9_Left_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Right_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_59_Left_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_53_Right_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_68_Left_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_62_Right_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_77_Left_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_71_Right_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_86_Left_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_80_Right_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTopModule_30 VGND VGND VPWR VPWR TopModule_30/HI Result[29] sky130_fd_sc_hd__conb_1
XFILLER_0_77_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_63_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_52_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTopModule_31 VGND VGND VPWR VPWR TopModule_31/HI Result[30] sky130_fd_sc_hd__conb_1
XTopModule_20 VGND VGND VPWR VPWR TopModule_20/HI Result[19] sky130_fd_sc_hd__conb_1
XFILLER_0_77_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_0_Left_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_39_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_368 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_81_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTopModule_21 VGND VGND VPWR VPWR TopModule_21/HI Result[20] sky130_fd_sc_hd__conb_1
XTopModule_10 VGND VGND VPWR VPWR TopModule_10/HI Result[9] sky130_fd_sc_hd__conb_1
XFILLER_0_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTopModule_32 VGND VGND VPWR VPWR TopModule_32/HI Result[31] sky130_fd_sc_hd__conb_1
XFILLER_0_77_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_19_Left_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_28_Left_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_37_Left_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_46_Left_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_55_Left_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_64_Left_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_73_Left_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_82_Left_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_81_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTopModule_22 VGND VGND VPWR VPWR TopModule_22/HI Result[21] sky130_fd_sc_hd__conb_1
XTopModule_11 VGND VGND VPWR VPWR TopModule_11/HI Result[10] sky130_fd_sc_hd__conb_1
XFILLER_0_77_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_69_Right_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_78_Right_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_68_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_87_Right_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_76_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_36_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTopModule_23 VGND VGND VPWR VPWR TopModule_23/HI Result[22] sky130_fd_sc_hd__conb_1
XFILLER_0_77_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTopModule_12 VGND VGND VPWR VPWR TopModule_12/HI Result[11] sky130_fd_sc_hd__conb_1
XFILLER_0_85_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_62_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_4_Left_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTopModule_24 VGND VGND VPWR VPWR TopModule_24/HI Result[23] sky130_fd_sc_hd__conb_1
XFILLER_0_77_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTopModule_13 VGND VGND VPWR VPWR TopModule_13/HI Result[12] sky130_fd_sc_hd__conb_1
XFILLER_0_85_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_39_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_86_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_15_Left_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_24_Left_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_33_Left_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_42_Left_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_51_Left_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_60_Left_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTopModule_25 VGND VGND VPWR VPWR TopModule_25/HI Result[24] sky130_fd_sc_hd__conb_1
XFILLER_0_85_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTopModule_14 VGND VGND VPWR VPWR TopModule_14/HI Result[13] sky130_fd_sc_hd__conb_1
XFILLER_0_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_94 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_47_Right_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_56_Right_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_65_Right_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_39_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_74_Right_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_89_Left_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_83_Right_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTopModule_26 VGND VGND VPWR VPWR TopModule_26/HI Result[25] sky130_fd_sc_hd__conb_1
XTopModule_15 VGND VGND VPWR VPWR TopModule_15/HI Result[14] sky130_fd_sc_hd__conb_1
XFILLER_0_73_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_8_Left_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_49_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_18_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTopModule_27 VGND VGND VPWR VPWR TopModule_27/HI Result[26] sky130_fd_sc_hd__conb_1
XTopModule_16 VGND VGND VPWR VPWR TopModule_16/HI Result[15] sky130_fd_sc_hd__conb_1
XFILLER_0_37_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Left_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Left_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_80_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_1_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTopModule_28 VGND VGND VPWR VPWR TopModule_28/HI Result[27] sky130_fd_sc_hd__conb_1
XTopModule_17 VGND VGND VPWR VPWR TopModule_17/HI Result[16] sky130_fd_sc_hd__conb_1
XFILLER_0_58_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_49_Left_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_43_Right_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_58_Left_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_52_Right_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_67_Left_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_61_Right_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_76_Left_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_70_Right_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_85_Left_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTopModule_29 VGND VGND VPWR VPWR TopModule_29/HI Result[28] sky130_fd_sc_hd__conb_1
XTopModule_18 VGND VGND VPWR VPWR TopModule_18/HI Result[17] sky130_fd_sc_hd__conb_1
XFILLER_0_58_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_30_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_86_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTopModule_19 VGND VGND VPWR VPWR TopModule_19/HI Result[18] sky130_fd_sc_hd__conb_1
XFILLER_0_37_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
.ends

