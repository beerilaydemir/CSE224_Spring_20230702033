magic
tech sky130A
magscale 1 2
timestamp 1748714431
<< nwell >>
rect 1066 2159 50086 51153
<< obsli1 >>
rect 1104 2159 50048 51153
<< obsm1 >>
rect 1104 2128 50218 51184
<< metal2 >>
rect 2226 52565 2282 53365
rect 5814 52565 5870 53365
rect 9402 52565 9458 53365
rect 12990 52565 13046 53365
rect 16578 52565 16634 53365
rect 20166 52565 20222 53365
rect 23754 52565 23810 53365
rect 27342 52565 27398 53365
rect 30930 52565 30986 53365
rect 34518 52565 34574 53365
rect 38106 52565 38162 53365
rect 41694 52565 41750 53365
rect 45282 52565 45338 53365
rect 48870 52565 48926 53365
<< obsm2 >>
rect 2338 52509 5758 52714
rect 5926 52509 9346 52714
rect 9514 52509 12934 52714
rect 13102 52509 16522 52714
rect 16690 52509 20110 52714
rect 20278 52509 23698 52714
rect 23866 52509 27286 52714
rect 27454 52509 30874 52714
rect 31042 52509 34462 52714
rect 34630 52509 38050 52714
rect 38218 52509 41638 52714
rect 41806 52509 45226 52714
rect 45394 52509 48814 52714
rect 48982 52509 50214 52714
rect 2282 2139 50214 52509
<< metal3 >>
rect 50421 49512 51221 49632
rect 50421 46792 51221 46912
rect 0 44072 800 44192
rect 50421 44072 51221 44192
rect 50421 41352 51221 41472
rect 50421 38632 51221 38752
rect 50421 35912 51221 36032
rect 50421 33192 51221 33312
rect 50421 30472 51221 30592
rect 50421 27752 51221 27872
rect 0 26392 800 26512
rect 50421 25032 51221 25152
rect 50421 22312 51221 22432
rect 50421 19592 51221 19712
rect 50421 16872 51221 16992
rect 50421 14152 51221 14272
rect 50421 11432 51221 11552
rect 0 8712 800 8832
rect 50421 8712 51221 8832
rect 50421 5992 51221 6112
rect 50421 3272 51221 3392
<< obsm3 >>
rect 4210 49712 50421 51169
rect 4210 49432 50341 49712
rect 4210 46992 50421 49432
rect 4210 46712 50341 46992
rect 4210 44272 50421 46712
rect 4210 43992 50341 44272
rect 4210 41552 50421 43992
rect 4210 41272 50341 41552
rect 4210 38832 50421 41272
rect 4210 38552 50341 38832
rect 4210 36112 50421 38552
rect 4210 35832 50341 36112
rect 4210 33392 50421 35832
rect 4210 33112 50341 33392
rect 4210 30672 50421 33112
rect 4210 30392 50341 30672
rect 4210 27952 50421 30392
rect 4210 27672 50341 27952
rect 4210 25232 50421 27672
rect 4210 24952 50341 25232
rect 4210 22512 50421 24952
rect 4210 22232 50341 22512
rect 4210 19792 50421 22232
rect 4210 19512 50341 19792
rect 4210 17072 50421 19512
rect 4210 16792 50341 17072
rect 4210 14352 50421 16792
rect 4210 14072 50341 14352
rect 4210 11632 50421 14072
rect 4210 11352 50341 11632
rect 4210 8912 50421 11352
rect 4210 8632 50341 8912
rect 4210 6192 50421 8632
rect 4210 5912 50341 6192
rect 4210 3472 50421 5912
rect 4210 3192 50341 3472
rect 4210 2143 50421 3192
<< metal4 >>
rect 4208 2128 4528 51184
rect 4868 2128 5188 51206
rect 5528 2128 5848 51184
rect 6188 2128 6508 51206
rect 6848 2128 7168 51184
rect 7508 2128 7828 51206
rect 8168 2128 8488 51184
rect 8828 2128 9148 51206
rect 9488 2128 9808 51184
rect 10148 2128 10468 51206
rect 10808 2128 11128 51184
rect 11468 2128 11788 51206
rect 12128 2128 12448 51184
rect 12788 2128 13108 51206
rect 13448 2128 13768 51184
rect 14108 2128 14428 51206
rect 14768 2128 15088 51184
rect 15428 2128 15748 51206
rect 16088 2128 16408 51184
rect 16748 2128 17068 51206
rect 17408 2128 17728 51184
rect 18068 2128 18388 51206
rect 18728 2128 19048 51184
rect 19388 2128 19708 51206
rect 20048 2128 20368 51184
rect 20708 2128 21028 51206
rect 21368 2128 21688 51184
rect 22028 2128 22348 51206
rect 22688 2128 23008 51184
rect 23348 2128 23668 51206
rect 24008 2128 24328 51184
rect 24668 2128 24988 51206
rect 25328 2128 25648 51184
rect 25988 2128 26308 51206
rect 26648 2128 26968 51184
rect 27308 2128 27628 51206
rect 27968 2128 28288 51184
rect 28628 2128 28948 51206
rect 29288 2128 29608 51184
rect 29948 2128 30268 51206
rect 30608 2128 30928 51184
rect 31268 2128 31588 51206
rect 31928 2128 32248 51184
rect 32588 2128 32908 51206
rect 33248 2128 33568 51184
rect 33908 2128 34228 51206
rect 34568 2128 34888 51184
rect 35228 2128 35548 51206
rect 35888 2128 36208 51184
rect 36548 2128 36868 51206
rect 37208 2128 37528 51184
rect 37868 2128 38188 51206
rect 38528 2128 38848 51184
rect 39188 2128 39508 51206
rect 39848 2128 40168 51184
rect 40508 2128 40828 51206
rect 41168 2128 41488 51184
rect 41828 2128 42148 51206
rect 42488 2128 42808 51184
rect 43148 2128 43468 51206
rect 43808 2128 44128 51184
rect 44468 2128 44788 51206
rect 45128 2128 45448 51184
rect 45788 2128 46108 51206
rect 46448 2128 46768 51184
rect 47108 2128 47428 51206
rect 47768 2128 48088 51184
rect 48428 2128 48748 51206
rect 49088 2128 49408 51184
rect 49748 2128 50068 51206
<< metal5 >>
rect 1056 50886 50096 51206
rect 1056 50226 50096 50546
rect 1056 49566 50096 49886
rect 1056 48906 50096 49226
rect 1056 48246 50096 48566
rect 1056 47586 50096 47906
rect 1056 46926 50096 47246
rect 1056 46266 50096 46586
rect 1056 45606 50096 45926
rect 1056 44946 50096 45266
rect 1056 44286 50096 44606
rect 1056 43626 50096 43946
rect 1056 42966 50096 43286
rect 1056 42306 50096 42626
rect 1056 41646 50096 41966
rect 1056 40986 50096 41306
rect 1056 40326 50096 40646
rect 1056 39666 50096 39986
rect 1056 39006 50096 39326
rect 1056 38346 50096 38666
rect 1056 37686 50096 38006
rect 1056 37026 50096 37346
rect 1056 36366 50096 36686
rect 1056 35706 50096 36026
rect 1056 35046 50096 35366
rect 1056 34386 50096 34706
rect 1056 33726 50096 34046
rect 1056 33066 50096 33386
rect 1056 32406 50096 32726
rect 1056 31746 50096 32066
rect 1056 31086 50096 31406
rect 1056 30426 50096 30746
rect 1056 29766 50096 30086
rect 1056 29106 50096 29426
rect 1056 28446 50096 28766
rect 1056 27786 50096 28106
rect 1056 27126 50096 27446
rect 1056 26466 50096 26786
rect 1056 25806 50096 26126
rect 1056 25146 50096 25466
rect 1056 24486 50096 24806
rect 1056 23826 50096 24146
rect 1056 23166 50096 23486
rect 1056 22506 50096 22826
rect 1056 21846 50096 22166
rect 1056 21186 50096 21506
rect 1056 20526 50096 20846
rect 1056 19866 50096 20186
rect 1056 19206 50096 19526
rect 1056 18546 50096 18866
rect 1056 17886 50096 18206
rect 1056 17226 50096 17546
rect 1056 16566 50096 16886
rect 1056 15906 50096 16226
rect 1056 15246 50096 15566
rect 1056 14586 50096 14906
rect 1056 13926 50096 14246
rect 1056 13266 50096 13586
rect 1056 12606 50096 12926
rect 1056 11946 50096 12266
rect 1056 11286 50096 11606
rect 1056 10626 50096 10946
rect 1056 9966 50096 10286
rect 1056 9306 50096 9626
rect 1056 8646 50096 8966
rect 1056 7986 50096 8306
rect 1056 7326 50096 7646
rect 1056 6666 50096 6986
rect 1056 6006 50096 6326
rect 1056 5346 50096 5666
<< labels >>
rlabel metal3 s 50421 3272 51221 3392 6 Result[0]
port 1 nsew signal output
rlabel metal3 s 50421 30472 51221 30592 6 Result[10]
port 2 nsew signal output
rlabel metal3 s 50421 33192 51221 33312 6 Result[11]
port 3 nsew signal output
rlabel metal3 s 50421 35912 51221 36032 6 Result[12]
port 4 nsew signal output
rlabel metal3 s 50421 38632 51221 38752 6 Result[13]
port 5 nsew signal output
rlabel metal3 s 50421 41352 51221 41472 6 Result[14]
port 6 nsew signal output
rlabel metal3 s 50421 44072 51221 44192 6 Result[15]
port 7 nsew signal output
rlabel metal3 s 50421 46792 51221 46912 6 Result[16]
port 8 nsew signal output
rlabel metal3 s 50421 49512 51221 49632 6 Result[17]
port 9 nsew signal output
rlabel metal2 s 2226 52565 2282 53365 6 Result[18]
port 10 nsew signal output
rlabel metal2 s 5814 52565 5870 53365 6 Result[19]
port 11 nsew signal output
rlabel metal3 s 50421 5992 51221 6112 6 Result[1]
port 12 nsew signal output
rlabel metal2 s 9402 52565 9458 53365 6 Result[20]
port 13 nsew signal output
rlabel metal2 s 12990 52565 13046 53365 6 Result[21]
port 14 nsew signal output
rlabel metal2 s 16578 52565 16634 53365 6 Result[22]
port 15 nsew signal output
rlabel metal2 s 20166 52565 20222 53365 6 Result[23]
port 16 nsew signal output
rlabel metal2 s 23754 52565 23810 53365 6 Result[24]
port 17 nsew signal output
rlabel metal2 s 27342 52565 27398 53365 6 Result[25]
port 18 nsew signal output
rlabel metal2 s 30930 52565 30986 53365 6 Result[26]
port 19 nsew signal output
rlabel metal2 s 34518 52565 34574 53365 6 Result[27]
port 20 nsew signal output
rlabel metal2 s 38106 52565 38162 53365 6 Result[28]
port 21 nsew signal output
rlabel metal2 s 41694 52565 41750 53365 6 Result[29]
port 22 nsew signal output
rlabel metal3 s 50421 8712 51221 8832 6 Result[2]
port 23 nsew signal output
rlabel metal2 s 45282 52565 45338 53365 6 Result[30]
port 24 nsew signal output
rlabel metal2 s 48870 52565 48926 53365 6 Result[31]
port 25 nsew signal output
rlabel metal3 s 50421 11432 51221 11552 6 Result[3]
port 26 nsew signal output
rlabel metal3 s 50421 14152 51221 14272 6 Result[4]
port 27 nsew signal output
rlabel metal3 s 50421 16872 51221 16992 6 Result[5]
port 28 nsew signal output
rlabel metal3 s 50421 19592 51221 19712 6 Result[6]
port 29 nsew signal output
rlabel metal3 s 50421 22312 51221 22432 6 Result[7]
port 30 nsew signal output
rlabel metal3 s 50421 25032 51221 25152 6 Result[8]
port 31 nsew signal output
rlabel metal3 s 50421 27752 51221 27872 6 Result[9]
port 32 nsew signal output
rlabel metal4 s 4868 2128 5188 51206 6 VGND
port 33 nsew ground bidirectional
rlabel metal4 s 6188 2128 6508 51206 6 VGND
port 33 nsew ground bidirectional
rlabel metal4 s 7508 2128 7828 51206 6 VGND
port 33 nsew ground bidirectional
rlabel metal4 s 8828 2128 9148 51206 6 VGND
port 33 nsew ground bidirectional
rlabel metal4 s 10148 2128 10468 51206 6 VGND
port 33 nsew ground bidirectional
rlabel metal4 s 11468 2128 11788 51206 6 VGND
port 33 nsew ground bidirectional
rlabel metal4 s 12788 2128 13108 51206 6 VGND
port 33 nsew ground bidirectional
rlabel metal4 s 14108 2128 14428 51206 6 VGND
port 33 nsew ground bidirectional
rlabel metal4 s 15428 2128 15748 51206 6 VGND
port 33 nsew ground bidirectional
rlabel metal4 s 16748 2128 17068 51206 6 VGND
port 33 nsew ground bidirectional
rlabel metal4 s 18068 2128 18388 51206 6 VGND
port 33 nsew ground bidirectional
rlabel metal4 s 19388 2128 19708 51206 6 VGND
port 33 nsew ground bidirectional
rlabel metal4 s 20708 2128 21028 51206 6 VGND
port 33 nsew ground bidirectional
rlabel metal4 s 22028 2128 22348 51206 6 VGND
port 33 nsew ground bidirectional
rlabel metal4 s 23348 2128 23668 51206 6 VGND
port 33 nsew ground bidirectional
rlabel metal4 s 24668 2128 24988 51206 6 VGND
port 33 nsew ground bidirectional
rlabel metal4 s 25988 2128 26308 51206 6 VGND
port 33 nsew ground bidirectional
rlabel metal4 s 27308 2128 27628 51206 6 VGND
port 33 nsew ground bidirectional
rlabel metal4 s 28628 2128 28948 51206 6 VGND
port 33 nsew ground bidirectional
rlabel metal4 s 29948 2128 30268 51206 6 VGND
port 33 nsew ground bidirectional
rlabel metal4 s 31268 2128 31588 51206 6 VGND
port 33 nsew ground bidirectional
rlabel metal4 s 32588 2128 32908 51206 6 VGND
port 33 nsew ground bidirectional
rlabel metal4 s 33908 2128 34228 51206 6 VGND
port 33 nsew ground bidirectional
rlabel metal4 s 35228 2128 35548 51206 6 VGND
port 33 nsew ground bidirectional
rlabel metal4 s 36548 2128 36868 51206 6 VGND
port 33 nsew ground bidirectional
rlabel metal4 s 37868 2128 38188 51206 6 VGND
port 33 nsew ground bidirectional
rlabel metal4 s 39188 2128 39508 51206 6 VGND
port 33 nsew ground bidirectional
rlabel metal4 s 40508 2128 40828 51206 6 VGND
port 33 nsew ground bidirectional
rlabel metal4 s 41828 2128 42148 51206 6 VGND
port 33 nsew ground bidirectional
rlabel metal4 s 43148 2128 43468 51206 6 VGND
port 33 nsew ground bidirectional
rlabel metal4 s 44468 2128 44788 51206 6 VGND
port 33 nsew ground bidirectional
rlabel metal4 s 45788 2128 46108 51206 6 VGND
port 33 nsew ground bidirectional
rlabel metal4 s 47108 2128 47428 51206 6 VGND
port 33 nsew ground bidirectional
rlabel metal4 s 48428 2128 48748 51206 6 VGND
port 33 nsew ground bidirectional
rlabel metal4 s 49748 2128 50068 51206 6 VGND
port 33 nsew ground bidirectional
rlabel metal5 s 1056 6006 50096 6326 6 VGND
port 33 nsew ground bidirectional
rlabel metal5 s 1056 7326 50096 7646 6 VGND
port 33 nsew ground bidirectional
rlabel metal5 s 1056 8646 50096 8966 6 VGND
port 33 nsew ground bidirectional
rlabel metal5 s 1056 9966 50096 10286 6 VGND
port 33 nsew ground bidirectional
rlabel metal5 s 1056 11286 50096 11606 6 VGND
port 33 nsew ground bidirectional
rlabel metal5 s 1056 12606 50096 12926 6 VGND
port 33 nsew ground bidirectional
rlabel metal5 s 1056 13926 50096 14246 6 VGND
port 33 nsew ground bidirectional
rlabel metal5 s 1056 15246 50096 15566 6 VGND
port 33 nsew ground bidirectional
rlabel metal5 s 1056 16566 50096 16886 6 VGND
port 33 nsew ground bidirectional
rlabel metal5 s 1056 17886 50096 18206 6 VGND
port 33 nsew ground bidirectional
rlabel metal5 s 1056 19206 50096 19526 6 VGND
port 33 nsew ground bidirectional
rlabel metal5 s 1056 20526 50096 20846 6 VGND
port 33 nsew ground bidirectional
rlabel metal5 s 1056 21846 50096 22166 6 VGND
port 33 nsew ground bidirectional
rlabel metal5 s 1056 23166 50096 23486 6 VGND
port 33 nsew ground bidirectional
rlabel metal5 s 1056 24486 50096 24806 6 VGND
port 33 nsew ground bidirectional
rlabel metal5 s 1056 25806 50096 26126 6 VGND
port 33 nsew ground bidirectional
rlabel metal5 s 1056 27126 50096 27446 6 VGND
port 33 nsew ground bidirectional
rlabel metal5 s 1056 28446 50096 28766 6 VGND
port 33 nsew ground bidirectional
rlabel metal5 s 1056 29766 50096 30086 6 VGND
port 33 nsew ground bidirectional
rlabel metal5 s 1056 31086 50096 31406 6 VGND
port 33 nsew ground bidirectional
rlabel metal5 s 1056 32406 50096 32726 6 VGND
port 33 nsew ground bidirectional
rlabel metal5 s 1056 33726 50096 34046 6 VGND
port 33 nsew ground bidirectional
rlabel metal5 s 1056 35046 50096 35366 6 VGND
port 33 nsew ground bidirectional
rlabel metal5 s 1056 36366 50096 36686 6 VGND
port 33 nsew ground bidirectional
rlabel metal5 s 1056 37686 50096 38006 6 VGND
port 33 nsew ground bidirectional
rlabel metal5 s 1056 39006 50096 39326 6 VGND
port 33 nsew ground bidirectional
rlabel metal5 s 1056 40326 50096 40646 6 VGND
port 33 nsew ground bidirectional
rlabel metal5 s 1056 41646 50096 41966 6 VGND
port 33 nsew ground bidirectional
rlabel metal5 s 1056 42966 50096 43286 6 VGND
port 33 nsew ground bidirectional
rlabel metal5 s 1056 44286 50096 44606 6 VGND
port 33 nsew ground bidirectional
rlabel metal5 s 1056 45606 50096 45926 6 VGND
port 33 nsew ground bidirectional
rlabel metal5 s 1056 46926 50096 47246 6 VGND
port 33 nsew ground bidirectional
rlabel metal5 s 1056 48246 50096 48566 6 VGND
port 33 nsew ground bidirectional
rlabel metal5 s 1056 49566 50096 49886 6 VGND
port 33 nsew ground bidirectional
rlabel metal5 s 1056 50886 50096 51206 6 VGND
port 33 nsew ground bidirectional
rlabel metal4 s 4208 2128 4528 51184 6 VPWR
port 34 nsew power bidirectional
rlabel metal4 s 5528 2128 5848 51184 6 VPWR
port 34 nsew power bidirectional
rlabel metal4 s 6848 2128 7168 51184 6 VPWR
port 34 nsew power bidirectional
rlabel metal4 s 8168 2128 8488 51184 6 VPWR
port 34 nsew power bidirectional
rlabel metal4 s 9488 2128 9808 51184 6 VPWR
port 34 nsew power bidirectional
rlabel metal4 s 10808 2128 11128 51184 6 VPWR
port 34 nsew power bidirectional
rlabel metal4 s 12128 2128 12448 51184 6 VPWR
port 34 nsew power bidirectional
rlabel metal4 s 13448 2128 13768 51184 6 VPWR
port 34 nsew power bidirectional
rlabel metal4 s 14768 2128 15088 51184 6 VPWR
port 34 nsew power bidirectional
rlabel metal4 s 16088 2128 16408 51184 6 VPWR
port 34 nsew power bidirectional
rlabel metal4 s 17408 2128 17728 51184 6 VPWR
port 34 nsew power bidirectional
rlabel metal4 s 18728 2128 19048 51184 6 VPWR
port 34 nsew power bidirectional
rlabel metal4 s 20048 2128 20368 51184 6 VPWR
port 34 nsew power bidirectional
rlabel metal4 s 21368 2128 21688 51184 6 VPWR
port 34 nsew power bidirectional
rlabel metal4 s 22688 2128 23008 51184 6 VPWR
port 34 nsew power bidirectional
rlabel metal4 s 24008 2128 24328 51184 6 VPWR
port 34 nsew power bidirectional
rlabel metal4 s 25328 2128 25648 51184 6 VPWR
port 34 nsew power bidirectional
rlabel metal4 s 26648 2128 26968 51184 6 VPWR
port 34 nsew power bidirectional
rlabel metal4 s 27968 2128 28288 51184 6 VPWR
port 34 nsew power bidirectional
rlabel metal4 s 29288 2128 29608 51184 6 VPWR
port 34 nsew power bidirectional
rlabel metal4 s 30608 2128 30928 51184 6 VPWR
port 34 nsew power bidirectional
rlabel metal4 s 31928 2128 32248 51184 6 VPWR
port 34 nsew power bidirectional
rlabel metal4 s 33248 2128 33568 51184 6 VPWR
port 34 nsew power bidirectional
rlabel metal4 s 34568 2128 34888 51184 6 VPWR
port 34 nsew power bidirectional
rlabel metal4 s 35888 2128 36208 51184 6 VPWR
port 34 nsew power bidirectional
rlabel metal4 s 37208 2128 37528 51184 6 VPWR
port 34 nsew power bidirectional
rlabel metal4 s 38528 2128 38848 51184 6 VPWR
port 34 nsew power bidirectional
rlabel metal4 s 39848 2128 40168 51184 6 VPWR
port 34 nsew power bidirectional
rlabel metal4 s 41168 2128 41488 51184 6 VPWR
port 34 nsew power bidirectional
rlabel metal4 s 42488 2128 42808 51184 6 VPWR
port 34 nsew power bidirectional
rlabel metal4 s 43808 2128 44128 51184 6 VPWR
port 34 nsew power bidirectional
rlabel metal4 s 45128 2128 45448 51184 6 VPWR
port 34 nsew power bidirectional
rlabel metal4 s 46448 2128 46768 51184 6 VPWR
port 34 nsew power bidirectional
rlabel metal4 s 47768 2128 48088 51184 6 VPWR
port 34 nsew power bidirectional
rlabel metal4 s 49088 2128 49408 51184 6 VPWR
port 34 nsew power bidirectional
rlabel metal5 s 1056 5346 50096 5666 6 VPWR
port 34 nsew power bidirectional
rlabel metal5 s 1056 6666 50096 6986 6 VPWR
port 34 nsew power bidirectional
rlabel metal5 s 1056 7986 50096 8306 6 VPWR
port 34 nsew power bidirectional
rlabel metal5 s 1056 9306 50096 9626 6 VPWR
port 34 nsew power bidirectional
rlabel metal5 s 1056 10626 50096 10946 6 VPWR
port 34 nsew power bidirectional
rlabel metal5 s 1056 11946 50096 12266 6 VPWR
port 34 nsew power bidirectional
rlabel metal5 s 1056 13266 50096 13586 6 VPWR
port 34 nsew power bidirectional
rlabel metal5 s 1056 14586 50096 14906 6 VPWR
port 34 nsew power bidirectional
rlabel metal5 s 1056 15906 50096 16226 6 VPWR
port 34 nsew power bidirectional
rlabel metal5 s 1056 17226 50096 17546 6 VPWR
port 34 nsew power bidirectional
rlabel metal5 s 1056 18546 50096 18866 6 VPWR
port 34 nsew power bidirectional
rlabel metal5 s 1056 19866 50096 20186 6 VPWR
port 34 nsew power bidirectional
rlabel metal5 s 1056 21186 50096 21506 6 VPWR
port 34 nsew power bidirectional
rlabel metal5 s 1056 22506 50096 22826 6 VPWR
port 34 nsew power bidirectional
rlabel metal5 s 1056 23826 50096 24146 6 VPWR
port 34 nsew power bidirectional
rlabel metal5 s 1056 25146 50096 25466 6 VPWR
port 34 nsew power bidirectional
rlabel metal5 s 1056 26466 50096 26786 6 VPWR
port 34 nsew power bidirectional
rlabel metal5 s 1056 27786 50096 28106 6 VPWR
port 34 nsew power bidirectional
rlabel metal5 s 1056 29106 50096 29426 6 VPWR
port 34 nsew power bidirectional
rlabel metal5 s 1056 30426 50096 30746 6 VPWR
port 34 nsew power bidirectional
rlabel metal5 s 1056 31746 50096 32066 6 VPWR
port 34 nsew power bidirectional
rlabel metal5 s 1056 33066 50096 33386 6 VPWR
port 34 nsew power bidirectional
rlabel metal5 s 1056 34386 50096 34706 6 VPWR
port 34 nsew power bidirectional
rlabel metal5 s 1056 35706 50096 36026 6 VPWR
port 34 nsew power bidirectional
rlabel metal5 s 1056 37026 50096 37346 6 VPWR
port 34 nsew power bidirectional
rlabel metal5 s 1056 38346 50096 38666 6 VPWR
port 34 nsew power bidirectional
rlabel metal5 s 1056 39666 50096 39986 6 VPWR
port 34 nsew power bidirectional
rlabel metal5 s 1056 40986 50096 41306 6 VPWR
port 34 nsew power bidirectional
rlabel metal5 s 1056 42306 50096 42626 6 VPWR
port 34 nsew power bidirectional
rlabel metal5 s 1056 43626 50096 43946 6 VPWR
port 34 nsew power bidirectional
rlabel metal5 s 1056 44946 50096 45266 6 VPWR
port 34 nsew power bidirectional
rlabel metal5 s 1056 46266 50096 46586 6 VPWR
port 34 nsew power bidirectional
rlabel metal5 s 1056 47586 50096 47906 6 VPWR
port 34 nsew power bidirectional
rlabel metal5 s 1056 48906 50096 49226 6 VPWR
port 34 nsew power bidirectional
rlabel metal5 s 1056 50226 50096 50546 6 VPWR
port 34 nsew power bidirectional
rlabel metal3 s 0 8712 800 8832 6 clk
port 35 nsew signal input
rlabel metal3 s 0 44072 800 44192 6 control
port 36 nsew signal input
rlabel metal3 s 0 26392 800 26512 6 reset
port 37 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 51221 53365
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 3808140
string GDS_FILE /openlane/designs/project5/runs/RUN_2025.05.31_18.00.03/results/signoff/TopModule.magic.gds
string GDS_START 23752
<< end >>

