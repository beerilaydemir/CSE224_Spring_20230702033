magic
tech sky130A
magscale 1 2
timestamp 1746885424
<< nwell >>
rect 1066 2159 18898 17425
<< obsli1 >>
rect 1104 2159 18860 17425
<< obsm1 >>
rect 106 484 19582 18828
<< metal2 >>
rect 1214 19200 1270 20000
rect 3698 19200 3754 20000
rect 6182 19200 6238 20000
rect 8666 19200 8722 20000
rect 11150 19200 11206 20000
rect 13634 19200 13690 20000
rect 16118 19200 16174 20000
rect 18602 19200 18658 20000
rect 3330 0 3386 800
rect 9954 0 10010 800
rect 16578 0 16634 800
<< obsm2 >>
rect 110 19144 1158 19200
rect 1326 19144 3642 19200
rect 3810 19144 6126 19200
rect 6294 19144 8610 19200
rect 8778 19144 11094 19200
rect 11262 19144 13578 19200
rect 13746 19144 16062 19200
rect 16230 19144 18546 19200
rect 18714 19144 19576 19200
rect 110 856 19576 19144
rect 110 439 3274 856
rect 3442 439 9898 856
rect 10066 439 16522 856
rect 16690 439 19576 856
<< metal3 >>
rect 0 18504 800 18624
rect 19200 18504 20000 18624
rect 0 16056 800 16176
rect 19200 16056 20000 16176
rect 0 13608 800 13728
rect 19200 13608 20000 13728
rect 0 11160 800 11280
rect 19200 11160 20000 11280
rect 0 8712 800 8832
rect 19200 8712 20000 8832
rect 0 6264 800 6384
rect 19200 6264 20000 6384
rect 0 3816 800 3936
rect 19200 3816 20000 3936
rect 0 1368 800 1488
rect 19200 1368 20000 1488
<< obsm3 >>
rect 105 18704 19450 18733
rect 880 18424 19120 18704
rect 105 16256 19450 18424
rect 880 15976 19120 16256
rect 105 13808 19450 15976
rect 880 13528 19120 13808
rect 105 11360 19450 13528
rect 880 11080 19120 11360
rect 105 8912 19450 11080
rect 880 8632 19120 8912
rect 105 6464 19450 8632
rect 880 6184 19120 6464
rect 105 4016 19450 6184
rect 880 3736 19120 4016
rect 105 1568 19450 3736
rect 880 1288 19120 1568
rect 105 443 19450 1288
<< metal4 >>
rect 1944 2128 2264 17456
rect 2604 2128 2924 17456
rect 6944 2128 7264 17456
rect 7604 2128 7924 17456
rect 11944 2128 12264 17456
rect 12604 2128 12924 17456
rect 16944 2128 17264 17456
rect 17604 2128 17924 17456
<< obsm4 >>
rect 795 17536 19530 18733
rect 795 2048 1864 17536
rect 2344 2048 2524 17536
rect 3004 2048 6864 17536
rect 7344 2048 7524 17536
rect 8004 2048 11864 17536
rect 12344 2048 12524 17536
rect 13004 2048 16864 17536
rect 17344 2048 17524 17536
rect 18004 2048 19530 17536
rect 795 443 19530 2048
<< metal5 >>
rect 1056 13676 18908 13996
rect 1056 13016 18908 13336
rect 1056 8676 18908 8996
rect 1056 8016 18908 8336
rect 1056 3676 18908 3996
rect 1056 3016 18908 3336
<< obsm5 >>
rect 852 14316 19572 16820
rect 19228 12696 19572 14316
rect 852 9316 19572 12696
rect 19228 7696 19572 9316
rect 852 4316 19572 7696
rect 19228 2696 19572 4316
rect 852 860 19572 2696
<< labels >>
rlabel metal3 s 0 18504 800 18624 6 A[0]
port 1 nsew signal input
rlabel metal3 s 0 16056 800 16176 6 A[1]
port 2 nsew signal input
rlabel metal3 s 0 13608 800 13728 6 A[2]
port 3 nsew signal input
rlabel metal3 s 0 11160 800 11280 6 A[3]
port 4 nsew signal input
rlabel metal3 s 0 8712 800 8832 6 A[4]
port 5 nsew signal input
rlabel metal3 s 0 6264 800 6384 6 A[5]
port 6 nsew signal input
rlabel metal3 s 0 3816 800 3936 6 A[6]
port 7 nsew signal input
rlabel metal3 s 0 1368 800 1488 6 A[7]
port 8 nsew signal input
rlabel metal2 s 18602 19200 18658 20000 6 B[0]
port 9 nsew signal input
rlabel metal2 s 16118 19200 16174 20000 6 B[1]
port 10 nsew signal input
rlabel metal2 s 13634 19200 13690 20000 6 B[2]
port 11 nsew signal input
rlabel metal2 s 11150 19200 11206 20000 6 B[3]
port 12 nsew signal input
rlabel metal2 s 8666 19200 8722 20000 6 B[4]
port 13 nsew signal input
rlabel metal2 s 6182 19200 6238 20000 6 B[5]
port 14 nsew signal input
rlabel metal2 s 3698 19200 3754 20000 6 B[6]
port 15 nsew signal input
rlabel metal2 s 1214 19200 1270 20000 6 B[7]
port 16 nsew signal input
rlabel metal4 s 2604 2128 2924 17456 6 VGND
port 17 nsew ground bidirectional
rlabel metal4 s 7604 2128 7924 17456 6 VGND
port 17 nsew ground bidirectional
rlabel metal4 s 12604 2128 12924 17456 6 VGND
port 17 nsew ground bidirectional
rlabel metal4 s 17604 2128 17924 17456 6 VGND
port 17 nsew ground bidirectional
rlabel metal5 s 1056 3676 18908 3996 6 VGND
port 17 nsew ground bidirectional
rlabel metal5 s 1056 8676 18908 8996 6 VGND
port 17 nsew ground bidirectional
rlabel metal5 s 1056 13676 18908 13996 6 VGND
port 17 nsew ground bidirectional
rlabel metal4 s 1944 2128 2264 17456 6 VPWR
port 18 nsew power bidirectional
rlabel metal4 s 6944 2128 7264 17456 6 VPWR
port 18 nsew power bidirectional
rlabel metal4 s 11944 2128 12264 17456 6 VPWR
port 18 nsew power bidirectional
rlabel metal4 s 16944 2128 17264 17456 6 VPWR
port 18 nsew power bidirectional
rlabel metal5 s 1056 3016 18908 3336 6 VPWR
port 18 nsew power bidirectional
rlabel metal5 s 1056 8016 18908 8336 6 VPWR
port 18 nsew power bidirectional
rlabel metal5 s 1056 13016 18908 13336 6 VPWR
port 18 nsew power bidirectional
rlabel metal2 s 16578 0 16634 800 6 opcode[0]
port 19 nsew signal input
rlabel metal2 s 9954 0 10010 800 6 opcode[1]
port 20 nsew signal input
rlabel metal2 s 3330 0 3386 800 6 opcode[2]
port 21 nsew signal input
rlabel metal3 s 19200 18504 20000 18624 6 out[0]
port 22 nsew signal output
rlabel metal3 s 19200 16056 20000 16176 6 out[1]
port 23 nsew signal output
rlabel metal3 s 19200 13608 20000 13728 6 out[2]
port 24 nsew signal output
rlabel metal3 s 19200 11160 20000 11280 6 out[3]
port 25 nsew signal output
rlabel metal3 s 19200 8712 20000 8832 6 out[4]
port 26 nsew signal output
rlabel metal3 s 19200 6264 20000 6384 6 out[5]
port 27 nsew signal output
rlabel metal3 s 19200 3816 20000 3936 6 out[6]
port 28 nsew signal output
rlabel metal3 s 19200 1368 20000 1488 6 out[7]
port 29 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 20000 20000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2065830
string GDS_FILE /openlane/designs/project2/runs/RUN_2025.05.10_13.53.11/results/signoff/alu.magic.gds
string GDS_START 601372
<< end >>

